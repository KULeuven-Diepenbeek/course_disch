    ...
    y(0) <= x(0) and x(1);
    y(1) <= x(2) and x(3);
    y(2) <= x(4) and x(5);
    y(3) <= x(6) and x(7);
    ...