my_shifted_vector(0) <= '0';
my_shifted_vector(1) <= '0';
my_shifted_vector(2) <= '0';
my_shifted_vector(3) <= my_vector(0);
my_shifted_vector(4) <= my_vector(1);
my_shifted_vector(5) <= my_vector(2);
my_shifted_vector(6) <= my_vector(3);
my_shifted_vector(7) <= my_vector(4);