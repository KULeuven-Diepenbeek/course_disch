
--------------------------------------------------------------------------------
-- KU Leuven - ESAT/COSIC - Emerging technologies, Systems & Security
--------------------------------------------------------------------------------
-- Module Name:     alu_tb - Behavioural
-- Project Name:    Testbench for alu
-- Description:     
--
-- Revision     Date       Author     Comments
-- v0.1         20240311   VlJo       Initial version
--
--------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
-- use IEEE.NUMERIC_STD.ALL;

entity alu_tb is
    generic(
        WIDTH : natural := 16
    );
end entity alu_tb;

architecture Behavioural of alu_tb is

    component alu is
        generic(
            WIDTH : natural := 16
        );
        port(
            X : IN STD_LOGIC_VECTOR(WIDTH-1 downto 0);
            Y : IN STD_LOGIC_VECTOR(WIDTH-1 downto 0);
            Z : OUT STD_LOGIC_VECTOR(WIDTH-1 downto 0);
            zx : IN STD_LOGIC;
            zy : IN STD_LOGIC;
            nx : IN STD_LOGIC;
            ny : IN STD_LOGIC;
            f : IN STD_LOGIC;
            no : IN STD_LOGIC;
            zr : OUT STD_LOGIC;
            ng : OUT STD_LOGIC
        );
    end component alu;

    signal X : STD_LOGIC_VECTOR(WIDTH-1 downto 0);
    signal Y : STD_LOGIC_VECTOR(WIDTH-1 downto 0);
    signal Z : STD_LOGIC_VECTOR(WIDTH-1 downto 0);
    signal zx : STD_LOGIC;
    signal zy : STD_LOGIC;
    signal nx : STD_LOGIC;
    signal ny : STD_LOGIC;
    signal f : STD_LOGIC;
    signal no : STD_LOGIC;
    signal zr : STD_LOGIC;
    signal ng : STD_LOGIC;

begin

    -------------------------------------------------------------------------------
    -- STIMULI
    -------------------------------------------------------------------------------
    PSTIM: process
    begin

        X <= x"0000";
        Y <= x"0000";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 10 ns;

        -- generate addition
        X <= x"c3fe";
        Y <= x"e4de";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3c02") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"7482";
        Y <= x"4bc7";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4082") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"aee5";
        Y <= x"068a";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"281d";
        Y <= x"02ad";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"fc60";
        Y <= x"feed";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"cf76";
        Y <= x"c71a";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"c719") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"b77c";
        Y <= x"a064";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"a064") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"8beb";
        Y <= x"8512";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7aee") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"8cb6";
        Y <= x"6e77";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"9189") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '1') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"c0e8";
        Y <= x"b315";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"b315") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"ff8b";
        Y <= x"8a84";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"757c") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"83ac";
        Y <= x"a4b8";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"5b48") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"f609";
        Y <= x"4b98";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4b97") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"d018";
        Y <= x"8228";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2fe7") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"12a6";
        Y <= x"97b9";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ed5a") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"10a3";
        Y <= x"bf97";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"bf96") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"6991";
        Y <= x"6299";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"06f8") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"0a32";
        Y <= x"4b6d";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4b7f") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '0') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"69c3";
        Y <= x"3986";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"c67a") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '1') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"4cb1";
        Y <= x"827d";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7d83") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"ac01";
        Y <= x"f887";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"fc87") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"70d2";
        Y <= x"a032";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"5fce") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"11a6";
        Y <= x"6ae3";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"f53f";
        Y <= x"7df0";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7df1") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"b732";
        Y <= x"b526";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"53e1";
        Y <= x"7818";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"5db7";
        Y <= x"4070";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4030") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"7061";
        Y <= x"d7e2";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"d7e1") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"80ad";
        Y <= x"ff81";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"007f") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"e1cb";
        Y <= x"323e";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"200a") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"ffc7";
        Y <= x"afbe";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"afbf") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"2dc9";
        Y <= x"4279";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"7042") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"4a7a";
        Y <= x"9f3f";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"60c0") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"e9f5";
        Y <= x"8751";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"160b") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"e8c0";
        Y <= x"5692";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"5693") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"655b";
        Y <= x"c270";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"5d15") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"98a9";
        Y <= x"dfdd";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2022") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"1a2f";
        Y <= x"16d4";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"16d5") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"0e3c";
        Y <= x"2d2e";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0c2c") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"e981";
        Y <= x"496e";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"496e") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"ba9c";
        Y <= x"495e";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b6a1") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"f1c5";
        Y <= x"9ab0";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f1c6") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"22e8";
        Y <= x"08ab";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"08ab") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"9964";
        Y <= x"1efa";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"eafd";
        Y <= x"b640";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"1502") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"331c";
        Y <= x"4ce0";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"6edc";
        Y <= x"6071";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"db98";
        Y <= x"1d3a";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"41a2") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"8b93";
        Y <= x"c994";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3e01") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"69ce";
        Y <= x"9271";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"69cf") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"a189";
        Y <= x"b01e";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"5e76") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"7326";
        Y <= x"7e7d";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"7e7c") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"c88f";
        Y <= x"bad7";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0db8") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"24ca";
        Y <= x"e443";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"e443") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"a9fb";
        Y <= x"0cf8";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"08f8") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"cee8";
        Y <= x"6448";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"cee7") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"011e";
        Y <= x"1fa2";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0102") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"46c4";
        Y <= x"0d61";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"c69d") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"0de5";
        Y <= x"6c7d";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"e207";
        Y <= x"304e";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"0254";
        Y <= x"98cb";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"fdac") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"6ff7";
        Y <= x"e4c7";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"6ff8") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"4af1";
        Y <= x"9544";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4af1") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"eb49";
        Y <= x"a41d";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a41e") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"a7b9";
        Y <= x"be8a";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"a7b8") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"c636";
        Y <= x"4e5e";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4e5f") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"2e95";
        Y <= x"6db6";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"b010";
        Y <= x"1ba9";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"4f01";
        Y <= x"84d5";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4f02") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"dfd0";
        Y <= x"ee7e";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2030") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"7709";
        Y <= x"d670";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"d670") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"4644";
        Y <= x"86f8";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"86f9") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"576c";
        Y <= x"9415";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"6beb") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"520c";
        Y <= x"9703";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"520b") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"466a";
        Y <= x"5fbb";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b995") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"ecb9";
        Y <= x"34d7";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"34d8") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"5660";
        Y <= x"83e3";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"f709";
        Y <= x"9411";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"08f7") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"26b7";
        Y <= x"291c";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"26b6") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"6f95";
        Y <= x"9767";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"9768") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"9d9a";
        Y <= x"bb9d";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"9998") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"97ea";
        Y <= x"e860";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"97eb") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"f697";
        Y <= x"bbc3";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"b25a") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"a47a";
        Y <= x"4613";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"5e67") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"dd52";
        Y <= x"3aac";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3aad") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"53ab";
        Y <= x"0b26";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f4d9") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"7049";
        Y <= x"cc84";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"5c3b") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"d044";
        Y <= x"6574";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"9530") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"1dcc";
        Y <= x"3779";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"1dcc") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"ab47";
        Y <= x"1499";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"54b9") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"2e31";
        Y <= x"012f";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2e30") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"8be0";
        Y <= x"d382";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2c7e") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"f165";
        Y <= x"8bc0";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"fbe5") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"05ee";
        Y <= x"06bc";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"5310";
        Y <= x"af53";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0263") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"01a9";
        Y <= x"68ed";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"fe56") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"b1c4";
        Y <= x"c078";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"d422";
        Y <= x"140b";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2bde") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"11c9";
        Y <= x"39d2";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"d7f7") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"34dc";
        Y <= x"c13c";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f618") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"c9ef";
        Y <= x"d200";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f7ef") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"f0d9";
        Y <= x"75b3";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f0d9") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"5697";
        Y <= x"0764";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"57f7") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '0') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"cd4e";
        Y <= x"3acd";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"32b1") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"da66";
        Y <= x"5efb";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"da65") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"f877";
        Y <= x"4b51";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ad26") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"e101";
        Y <= x"d68a";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0a77") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"3e05";
        Y <= x"c2f8";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"6579";
        Y <= x"d88b";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"9a87") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"2609";
        Y <= x"8bfb";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"260a") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"34e8";
        Y <= x"b799";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4866") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"1178";
        Y <= x"28a0";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"28a0") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"1688";
        Y <= x"706c";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"61a0";
        Y <= x"1569";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"619f") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"64a8";
        Y <= x"d517";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"d516") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"1040";
        Y <= x"4d21";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b2de") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"a8b9";
        Y <= x"4b03";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4b03") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"fd3f";
        Y <= x"7eaf";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7eb0") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"048d";
        Y <= x"0348";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0008") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"07bc";
        Y <= x"0173";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f9b7") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"f0ae";
        Y <= x"e608";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f0af") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"12fd";
        Y <= x"eedf";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"eee0") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"5f61";
        Y <= x"746f";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a09e") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"5b42";
        Y <= x"34d4";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a4bd") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"1014";
        Y <= x"64ef";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"5c9a";
        Y <= x"a3ca";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a3cb") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"c414";
        Y <= x"8407";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"c414") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"35aa";
        Y <= x"8fe5";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"35ab") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"1006";
        Y <= x"f94d";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"16b9") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"994e";
        Y <= x"4c89";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"994f") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"3a4e";
        Y <= x"e139";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e13a") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"964e";
        Y <= x"b0fc";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"474a") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"0c45";
        Y <= x"bc04";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0c44") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"8acc";
        Y <= x"e272";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"8240") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"2d2c";
        Y <= x"c2fb";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"0ae7";
        Y <= x"5036";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"5b1d") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"fa6b";
        Y <= x"2c2e";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"fe6f") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"c441";
        Y <= x"cf27";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"c441") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"84da";
        Y <= x"a485";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"5b7b") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"854b";
        Y <= x"531c";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"ab5a";
        Y <= x"7a68";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"54a5") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"0f11";
        Y <= x"e3b5";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"efb5") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"3bf7";
        Y <= x"9571";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3bf8") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"66b7";
        Y <= x"0033";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0033") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"86d5";
        Y <= x"df07";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"8605") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"4a65";
        Y <= x"d435";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"d435") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"bd56";
        Y <= x"7561";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"fd77") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"16c2";
        Y <= x"07f8";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"07f7") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"42ee";
        Y <= x"5556";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"42ee") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"5753";
        Y <= x"4696";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4697") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"22b3";
        Y <= x"9704";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"b9b7") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"716a";
        Y <= x"94f3";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"94f4") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"00d2";
        Y <= x"f824";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f752") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"3937";
        Y <= x"ce0d";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"c6c9") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"e965";
        Y <= x"afd5";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"993a") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"e9d7";
        Y <= x"dd4d";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"1628") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"9c6c";
        Y <= x"f4c5";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f4c4") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"89a1";
        Y <= x"6795";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"efb5") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"b9a0";
        Y <= x"b16a";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0836") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"7c8b";
        Y <= x"0f42";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f0bd") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"46cf";
        Y <= x"1e61";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"7977";
        Y <= x"7f1f";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"8689") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"6261";
        Y <= x"21e8";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"f107";
        Y <= x"dde5";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"d105") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"5804";
        Y <= x"2942";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2943") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"f606";
        Y <= x"a9e4";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f607") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"9ffc";
        Y <= x"703e";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"703e") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"943f";
        Y <= x"22ac";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"b6eb") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"7443";
        Y <= x"749f";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"2313";
        Y <= x"a36a";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2302") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"c1e2";
        Y <= x"8923";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"c1e2") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"308b";
        Y <= x"eea4";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"cf75") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"8c14";
        Y <= x"bbbb";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"8810") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"5549";
        Y <= x"577a";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"5779") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"cb93";
        Y <= x"6cd3";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a140") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"5c06";
        Y <= x"25fd";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7dff") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '0') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"4cba";
        Y <= x"7adc";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"7adb") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"5a57";
        Y <= x"44a7";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"5a57") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"6c81";
        Y <= x"7691";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"8a15";
        Y <= x"d9aa";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"dbbf") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"9654";
        Y <= x"caeb";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"caec") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"6e4b";
        Y <= x"47fa";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"47f9") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"45fe";
        Y <= x"fa60";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"8c79";
        Y <= x"4a1f";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"d1dc";
        Y <= x"4382";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"71a6") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"77bc";
        Y <= x"c9b9";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ae03") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"b71d";
        Y <= x"c5c1";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"48e3") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"681a";
        Y <= x"37d0";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"d7e6";
        Y <= x"8b89";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"281a") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"7f5d";
        Y <= x"4998";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"7f5c") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"0f23";
        Y <= x"20d9";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ee4a") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"c506";
        Y <= x"3ab6";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"c54a") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '1') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"7395";
        Y <= x"77ed";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"77fd") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '0') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"b581";
        Y <= x"efc8";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"a549") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"7c22";
        Y <= x"b6c4";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"493c") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"45d5";
        Y <= x"732a";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"45d6") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"72f2";
        Y <= x"301e";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"d12c";
        Y <= x"2c95";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0004") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"afbe";
        Y <= x"5eb3";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0eb2") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"1aab";
        Y <= x"ad72";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"1aab") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"17d6";
        Y <= x"f8aa";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"79d3";
        Y <= x"570b";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a8f5") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '1') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"dae8";
        Y <= x"dcc7";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"dcc7") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"f06f";
        Y <= x"c624";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0f90") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"9d71";
        Y <= x"5947";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"b2f1";
        Y <= x"ccf7";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e5fa") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"abcc";
        Y <= x"90b9";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"5f47";
        Y <= x"0585";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0585") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"5232";
        Y <= x"974a";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"974b") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"9d06";
        Y <= x"e87d";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"1783") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"40ee";
        Y <= x"ed24";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ac36") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"7833";
        Y <= x"1a0f";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e5f0") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"f574";
        Y <= x"02dd";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f574") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"af24";
        Y <= x"f423";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f424") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"1848";
        Y <= x"ac34";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"53cb") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"2a61";
        Y <= x"06f8";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2a61") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"35a3";
        Y <= x"ac67";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ac68") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"69a6";
        Y <= x"3b0f";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"3b0f") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"3f7c";
        Y <= x"c868";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"3f7b") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"78ac";
        Y <= x"f174";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"78ab") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"f3fe";
        Y <= x"37a0";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f7fe") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"ec28";
        Y <= x"728a";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"8c38";
        Y <= x"954c";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"954c") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"5198";
        Y <= x"b6a0";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"5197") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"4d92";
        Y <= x"bddd";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"8fb5") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"0988";
        Y <= x"e877";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0989") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"c201";
        Y <= x"fa62";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"c202") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"7035";
        Y <= x"8abb";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0031") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"f842";
        Y <= x"45ff";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f842") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"4834";
        Y <= x"e7fd";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e7fe") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"5110";
        Y <= x"43f7";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0d19") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"63f3";
        Y <= x"3289";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"9c0c") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"05d4";
        Y <= x"b050";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"05d4") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"3ef7";
        Y <= x"a72f";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3ef8") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"39a2";
        Y <= x"b0cc";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"39a3") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"8111";
        Y <= x"b570";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"cba1") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"8ffe";
        Y <= x"4a34";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4a33") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"356c";
        Y <= x"a82b";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"356d") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"f820";
        Y <= x"c2ae";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"07e0") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"d8ba";
        Y <= x"0a25";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"e2df") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"48f3";
        Y <= x"80d7";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"48f4") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"9337";
        Y <= x"1989";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"acc0") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"179c";
        Y <= x"cc60";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b4c4") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"91c8";
        Y <= x"791b";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"6e37") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"2029";
        Y <= x"6b8c";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"6bad") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '0') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"0128";
        Y <= x"0148";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0147") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"50e0";
        Y <= x"b541";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4abf") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"eea4";
        Y <= x"07e0";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"115b") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"32f4";
        Y <= x"91cf";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"32f4") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"6a18";
        Y <= x"1707";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"1707") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"6991";
        Y <= x"2fa4";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"c613") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"5588";
        Y <= x"ef8a";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"c915";
        Y <= x"f66a";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"c000") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"c276";
        Y <= x"d7f4";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"280b") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"b191";
        Y <= x"656e";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"656d") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"1b62";
        Y <= x"eee4";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"ba4d";
        Y <= x"a9e3";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"45b2") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"b706";
        Y <= x"5e06";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a700") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"f0c4";
        Y <= x"9f1e";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"9f1e") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"769e";
        Y <= x"125b";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"769f") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"0bac";
        Y <= x"8fda";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7026") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"51c0";
        Y <= x"d4d8";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"c624";
        Y <= x"5ef2";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"def6") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"8096";
        Y <= x"f15d";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"d898";
        Y <= x"c219";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"da99") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"8833";
        Y <= x"3d7e";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"77cc") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"946b";
        Y <= x"aab5";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"aab4") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"6513";
        Y <= x"ea78";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"1587") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"ed1b";
        Y <= x"526d";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"12e5") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"69fd";
        Y <= x"7db4";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"9602") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"6078";
        Y <= x"f1dd";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f1dd") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"fcc7";
        Y <= x"f288";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f288") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"0cf9";
        Y <= x"a41b";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"b114") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"d7b2";
        Y <= x"b48f";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"284d") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"b63c";
        Y <= x"b383";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"b382") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"4a56";
        Y <= x"8d90";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"8d8f") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"e1d7";
        Y <= x"ee10";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"11f0") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"ac2b";
        Y <= x"8829";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2402") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"c39a";
        Y <= x"50a6";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"af5a") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '1') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"339b";
        Y <= x"ad51";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"52ae") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"5490";
        Y <= x"6b73";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"fd7a";
        Y <= x"6c4f";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"fd7a") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"b81b";
        Y <= x"dde9";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"25ce") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"02ed";
        Y <= x"7f69";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"02ee") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"801b";
        Y <= x"1ebb";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"381f";
        Y <= x"c7b9";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"381f") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"7ecc";
        Y <= x"daf5";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"383d";
        Y <= x"b6cd";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"300d") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"eb5c";
        Y <= x"42b8";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"b5ba";
        Y <= x"ec6b";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b5bb") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"0150";
        Y <= x"5484";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"feaf") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"ae4e";
        Y <= x"a490";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f642") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"f379";
        Y <= x"b6ac";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"aa25") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"12f3";
        Y <= x"db7c";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"12f4") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"5c0e";
        Y <= x"e252";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a3f1") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"deb8";
        Y <= x"28a8";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"982c";
        Y <= x"d97b";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"d97b") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"0083";
        Y <= x"09a0";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ff7d") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"75e8";
        Y <= x"a0c3";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"def2";
        Y <= x"d3f6";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"655f";
        Y <= x"3ec8";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"6560") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"657c";
        Y <= x"8071";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"e5ed") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"0f97";
        Y <= x"3cdd";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f069") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"e551";
        Y <= x"2e5f";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"d1a1") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '1') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"396d";
        Y <= x"1326";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"396c") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"fd39";
        Y <= x"b08d";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"02c6") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"08a9";
        Y <= x"039a";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0088") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"c643";
        Y <= x"f916";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f916") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"d206";
        Y <= x"fa7d";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"fa7f") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"932a";
        Y <= x"d9a1";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"d9a0") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"95a3";
        Y <= x"fcc7";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"6a5c") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"bbba";
        Y <= x"8538";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"951d";
        Y <= x"d237";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"c2e6") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"d011";
        Y <= x"a23a";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"1f10";
        Y <= x"822d";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7dd2") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"368f";
        Y <= x"0443";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"a07c";
        Y <= x"69d7";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"ec6b";
        Y <= x"393b";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"1395") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"d3bd";
        Y <= x"cc92";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"336d") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"a50e";
        Y <= x"5988";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"c732";
        Y <= x"ac73";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e541") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"c59a";
        Y <= x"8174";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"c59a") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"5be1";
        Y <= x"cb48";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"34b8") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"375d";
        Y <= x"e93e";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e93f") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"3ebc";
        Y <= x"b64a";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"3ebc") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"71b6";
        Y <= x"002e";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"de4c";
        Y <= x"5cbc";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"21b4") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"34cc";
        Y <= x"7121";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3c55") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"42cb";
        Y <= x"b6f8";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"b736";
        Y <= x"56c5";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a93b") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '1') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"552d";
        Y <= x"5f40";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"45b5";
        Y <= x"3dde";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"45b4") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"1a4c";
        Y <= x"bb2b";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"5f21") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"3145";
        Y <= x"8943";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"af19";
        Y <= x"8af9";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7506") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"0115";
        Y <= x"6db4";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"feea") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"4b8f";
        Y <= x"71b5";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7bbf") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '0') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"18fc";
        Y <= x"e305";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"09a4";
        Y <= x"aed3";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a52f") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"7fa6";
        Y <= x"adce";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"adce") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"3c0d";
        Y <= x"c89d";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"3c0d") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"a7ac";
        Y <= x"c1bf";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"5854") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"4459";
        Y <= x"abfd";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4458") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"7fd0";
        Y <= x"7f05";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7fd1") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"07b1";
        Y <= x"0962";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f69d") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"fe22";
        Y <= x"c5b3";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"01de") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"b842";
        Y <= x"7a62";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"47bd") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"4368";
        Y <= x"3e69";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4369") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"5e25";
        Y <= x"b30a";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"4d2d";
        Y <= x"675f";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"b48c") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"6280";
        Y <= x"ac10";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2000") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"4d1f";
        Y <= x"ef7a";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4d1f") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"f28e";
        Y <= x"0109";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"fef6") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"3812";
        Y <= x"59e5";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a61a") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"9b42";
        Y <= x"49c7";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0942") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"f76b";
        Y <= x"cba7";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0895") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"a22c";
        Y <= x"2ba6";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"d459") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"5972";
        Y <= x"f586";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a68d") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"887a";
        Y <= x"8a87";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"8a88") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"348d";
        Y <= x"6c04";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"6c03") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"b883";
        Y <= x"a2a6";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"a082") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"8855";
        Y <= x"8d7a";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"8850") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"d45e";
        Y <= x"96ff";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"182c";
        Y <= x"0fb1";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"182d") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"7a22";
        Y <= x"8813";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"77ec") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"d94f";
        Y <= x"f028";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"d2de";
        Y <= x"f859";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"fadf") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"2fcc";
        Y <= x"c55d";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f529") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"4bde";
        Y <= x"02ab";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4bdd") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"c915";
        Y <= x"278d";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"36eb") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"d77e";
        Y <= x"3a27";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"ba8c";
        Y <= x"7766";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"bcda") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"8c69";
        Y <= x"7f87";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7f88") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"63a0";
        Y <= x"9aad";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"6553") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"a300";
        Y <= x"3388";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"cc77") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"ed2b";
        Y <= x"ea5b";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"15a4") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"496e";
        Y <= x"b5c9";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"fdef";
        Y <= x"79e2";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"79e1") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"1437";
        Y <= x"6326";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4eef") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"b4c5";
        Y <= x"cf1d";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"83e2") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"fa42";
        Y <= x"5707";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"05be") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"524e";
        Y <= x"bb46";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"44ba") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"639c";
        Y <= x"e3da";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"639d") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"76c8";
        Y <= x"ee4c";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ee4d") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"8bba";
        Y <= x"9d80";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"8980") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"22bf";
        Y <= x"a8d5";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"a8d4") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"fd50";
        Y <= x"8979";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"8c29") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"d6c9";
        Y <= x"4e6b";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b195") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '1') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"76d6";
        Y <= x"fc04";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"8929") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"288b";
        Y <= x"a8ed";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"d774") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"815d";
        Y <= x"50db";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"815e") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"01e8";
        Y <= x"7a44";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"7a43") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"7525";
        Y <= x"73db";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"014a") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"eecf";
        Y <= x"42a8";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"8d2a";
        Y <= x"f6e1";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ffeb") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"7b78";
        Y <= x"bcae";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"bcaf") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"2128";
        Y <= x"3abb";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2028") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"cdf0";
        Y <= x"c3a3";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"cdef") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"114d";
        Y <= x"3235";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"cdcb") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '1') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"052d";
        Y <= x"4638";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"d44b";
        Y <= x"5e23";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2bb5") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"babe";
        Y <= x"ba9e";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"babf") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"577a";
        Y <= x"592f";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"512a") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"a9a4";
        Y <= x"2cb2";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"28a0") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"35da";
        Y <= x"78fc";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4322") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"159e";
        Y <= x"a6db";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"4e7c";
        Y <= x"8050";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ce7c") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"b510";
        Y <= x"3728";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"8218") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"38ba";
        Y <= x"ed84";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2880") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"22e2";
        Y <= x"a962";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"a961") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"8492";
        Y <= x"6ef5";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f387") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"60b4";
        Y <= x"1213";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"60b4") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"2c0d";
        Y <= x"778a";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"8876") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '1') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"f004";
        Y <= x"008c";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f004") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"98d2";
        Y <= x"699c";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"98d3") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"2676";
        Y <= x"1964";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"dbc3";
        Y <= x"f99b";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f99c") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"45ef";
        Y <= x"a056";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a057") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"1cbe";
        Y <= x"94a0";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"881e") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"d831";
        Y <= x"a413";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"27cf") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"5168";
        Y <= x"b47d";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4b82") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"7631";
        Y <= x"5641";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"9532";
        Y <= x"cd73";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"8532") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"1fa6";
        Y <= x"8277";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"62d1") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"afb1";
        Y <= x"b78e";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"07dd") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"bd53";
        Y <= x"9052";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"9052") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"d3b7";
        Y <= x"1b9d";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"1b9d") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"dd77";
        Y <= x"0267";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"dfde") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"24c1";
        Y <= x"783e";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"24c0") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"e158";
        Y <= x"ce55";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e159") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"ebf0";
        Y <= x"4a8e";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b571") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"53ea";
        Y <= x"2ba4";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ac15") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"cac7";
        Y <= x"1af5";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"502e") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"ae72";
        Y <= x"9642";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ae71") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"4f98";
        Y <= x"2f31";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0f10") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"d9e6";
        Y <= x"367d";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"ca05";
        Y <= x"1ca6";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e35a") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '1') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"549b";
        Y <= x"383e";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"8e1c";
        Y <= x"f49f";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"71e3") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"e0fa";
        Y <= x"e944";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"16bb") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"56a4";
        Y <= x"c120";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"3af5";
        Y <= x"bd84";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"3884") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"6578";
        Y <= x"5f89";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"5e6d";
        Y <= x"44a9";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"19c4") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"dea1";
        Y <= x"5579";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"dea1") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"81d2";
        Y <= x"a9e8";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"81c0") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"e932";
        Y <= x"dd83";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"16cd") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"004d";
        Y <= x"9db5";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"9e02") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"6f09";
        Y <= x"45d5";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"6fdd") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '0') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"70c4";
        Y <= x"f216";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"70c4") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"f223";
        Y <= x"fbe8";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"fbe9") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"cdd6";
        Y <= x"0956";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"cdd6") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"3235";
        Y <= x"a321";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"a320") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"de03";
        Y <= x"f0f1";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f0f1") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"2c1a";
        Y <= x"33a3";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"2398";
        Y <= x"ac4c";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"afdc") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"ee6d";
        Y <= x"c073";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"1192") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"d1a7";
        Y <= x"702f";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"9e88") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"59a0";
        Y <= x"6c20";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"6c1f") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"d07c";
        Y <= x"e9ee";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"1611") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"3ac6";
        Y <= x"37d2";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"f374";
        Y <= x"5630";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f373") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"85fe";
        Y <= x"e23a";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"1dc5") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"a3d6";
        Y <= x"edca";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"a1c2") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"1994";
        Y <= x"c0ca";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3f36") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"9451";
        Y <= x"2967";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"9452") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"c7d0";
        Y <= x"5a16";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"5a15") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"72d8";
        Y <= x"6685";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"6684") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"3d8e";
        Y <= x"66c7";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3d8f") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"a2f4";
        Y <= x"e17d";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e17e") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"a562";
        Y <= x"8bae";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a563") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"7d69";
        Y <= x"9ce6";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"8297") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"a818";
        Y <= x"c303";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"57e8") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"732c";
        Y <= x"3063";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"8cd4") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"5d02";
        Y <= x"182b";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"5d02") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"559b";
        Y <= x"2d72";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2d71") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"fab4";
        Y <= x"3d85";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"c27a") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"89b3";
        Y <= x"f863";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"764c") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"d81e";
        Y <= x"a7a8";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"8008") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"f84b";
        Y <= x"3b3e";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"c4c1") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"a235";
        Y <= x"e06e";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a236") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"11c8";
        Y <= x"f355";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"1e73") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"49c6";
        Y <= x"987e";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"8d9a";
        Y <= x"a921";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"fb10";
        Y <= x"ab88";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"9f1d";
        Y <= x"ed1e";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"9c6c";
        Y <= x"b05c";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"2382";
        Y <= x"1d4c";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3fce") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '0') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"b75e";
        Y <= x"12d0";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"48a1") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"ab2d";
        Y <= x"409a";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"bf66") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '1') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"fd36";
        Y <= x"6215";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"6014") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"eeb2";
        Y <= x"aa32";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"eeb1") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"f4e1";
        Y <= x"a5d0";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"5b98";
        Y <= x"30e2";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"30e1") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"7ebc";
        Y <= x"8ff5";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"8ff6") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"6621";
        Y <= x"4be5";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4be5") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"3ebb";
        Y <= x"62a8";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"c145") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"1060";
        Y <= x"f7fd";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"3bc8";
        Y <= x"74fa";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"3bc8") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"219a";
        Y <= x"b3ad";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"de65") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"50b5";
        Y <= x"1357";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3d5e") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"f982";
        Y <= x"567c";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a306") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"54d7";
        Y <= x"bb9a";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4465") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"a28f";
        Y <= x"a93f";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"5d70") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"9f21";
        Y <= x"fc0e";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"60df") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"788e";
        Y <= x"a270";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"7be1";
        Y <= x"92af";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"92af") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"bf87";
        Y <= x"6ce7";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"52a0") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"c2f6";
        Y <= x"9a8d";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3d0a") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"4853";
        Y <= x"4031";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0822") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"35dc";
        Y <= x"1be5";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"35db") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"3d94";
        Y <= x"832e";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3d95") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"29ef";
        Y <= x"ec63";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"1652") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"ed2b";
        Y <= x"59b9";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"e00e";
        Y <= x"ae86";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"4a10";
        Y <= x"e4da";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"563b";
        Y <= x"e246";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"73f5") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"6e8e";
        Y <= x"bc76";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"6e8d") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"e044";
        Y <= x"2a53";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"1fbb") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"44fe";
        Y <= x"29e2";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"d61d") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"6e62";
        Y <= x"0166";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"6fc8") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"ff2b";
        Y <= x"0d34";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0c5f") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"cfbe";
        Y <= x"4cc0";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"fe43";
        Y <= x"19f4";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"1a63";
        Y <= x"a725";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"58db") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"c2dc";
        Y <= x"e431";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"e431") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"bfdc";
        Y <= x"9a96";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"0054";
        Y <= x"9d27";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"bf85";
        Y <= x"e466";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"24e1") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"f7ae";
        Y <= x"169a";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e114") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"4239";
        Y <= x"a0ea";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4238") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"2344";
        Y <= x"613a";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"9ec5") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"5f00";
        Y <= x"0116";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0100") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"fbac";
        Y <= x"c05e";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"fbab") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"7ff7";
        Y <= x"bec0";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4140") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"a4c0";
        Y <= x"e18f";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"a080") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"b243";
        Y <= x"c3a4";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3c5b") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"369e";
        Y <= x"5870";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"369e") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"fad3";
        Y <= x"36b4";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"00b9";
        Y <= x"e489";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"3aff";
        Y <= x"c5a3";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"00a2") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"46cf";
        Y <= x"a7a1";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0681") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"3247";
        Y <= x"4d1c";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"3246") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"b468";
        Y <= x"5cb8";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b469") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"00c1";
        Y <= x"4577";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ba89") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '1') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"5fee";
        Y <= x"4d94";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4d94") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"3ddd";
        Y <= x"22c2";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"e051";
        Y <= x"a2b9";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"d482";
        Y <= x"8a8b";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"650a";
        Y <= x"bf58";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"5a4e") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"ca98";
        Y <= x"d792";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"d791") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"fcd8";
        Y <= x"a40a";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"a408") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"7adc";
        Y <= x"add3";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"f8a9";
        Y <= x"f7a1";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f8a8") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"84f0";
        Y <= x"f435";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"84ef") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"4782";
        Y <= x"ef1f";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b87d") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"cdcc";
        Y <= x"efa3";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"efa2") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"9ced";
        Y <= x"a689";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"a689") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"7091";
        Y <= x"95c3";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"dace") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"6d4a";
        Y <= x"b1b4";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"b1b4") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"2159";
        Y <= x"c8ba";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"35e2";
        Y <= x"1d3f";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"1522") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"5123";
        Y <= x"b51a";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"aedd") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"685f";
        Y <= x"ab8f";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"69c2";
        Y <= x"c1ca";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"69c2") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"9f52";
        Y <= x"875e";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"9f51") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"587f";
        Y <= x"c051";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a780") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"aeb2";
        Y <= x"dcd1";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"6340";
        Y <= x"d90a";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"cc4a";
        Y <= x"849a";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"849b") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"e9c3";
        Y <= x"c060";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"e9c2") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"0872";
        Y <= x"6c8e";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0871") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"d96a";
        Y <= x"b6f4";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2695") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"7eb4";
        Y <= x"d2a1";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"814c") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"3040";
        Y <= x"31be";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"1ca5";
        Y <= x"16d5";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"337a") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"fdab";
        Y <= x"02f1";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"fdaa") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"60e1";
        Y <= x"1fd1";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"9f1f") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"c756";
        Y <= x"b3cd";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"38a9") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"f42c";
        Y <= x"ae94";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"516b") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"e50d";
        Y <= x"9d18";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"62e8") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"9243";
        Y <= x"96fc";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"6903") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"948f";
        Y <= x"1533";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"7db0";
        Y <= x"2db4";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"1203";
        Y <= x"233a";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"1203") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"09ff";
        Y <= x"09be";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ffbf") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"1c6c";
        Y <= x"576a";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e393") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"14a0";
        Y <= x"3154";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"14a0") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"a247";
        Y <= x"88b8";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7748") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"2963";
        Y <= x"e0cf";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2963") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"3bff";
        Y <= x"bb58";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"5aab";
        Y <= x"d84d";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a555") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"9c9c";
        Y <= x"e303";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"6363") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"25ad";
        Y <= x"5fd1";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"572a";
        Y <= x"d320";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"572b") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"ddb5";
        Y <= x"a65d";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"224b") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"ea4c";
        Y <= x"7a10";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"703c") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"e3bb";
        Y <= x"0b85";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ef40") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"0e19";
        Y <= x"5d91";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4f78") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"7397";
        Y <= x"ce70";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4210") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"34d4";
        Y <= x"c6b6";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"fb8a") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"55b1";
        Y <= x"8d42";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"7211";
        Y <= x"a31e";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"cde6";
        Y <= x"4af8";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4af8") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"0c94";
        Y <= x"c4ec";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3b13") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"e4d7";
        Y <= x"208d";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"208d") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"6014";
        Y <= x"acb7";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"6013") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"4090";
        Y <= x"38e7";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4091") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"6df8";
        Y <= x"c65b";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"9208") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"c20d";
        Y <= x"402f";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"023c") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"c872";
        Y <= x"2d72";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f5e4") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"1ff0";
        Y <= x"9891";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e00f") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"c34d";
        Y <= x"35ae";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"35af") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"7e83";
        Y <= x"c6e3";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"391d") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"f0a1";
        Y <= x"ea76";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f0a1") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"a8b1";
        Y <= x"c2ff";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"6bb0") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"5236";
        Y <= x"3041";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"3041") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"fc57";
        Y <= x"42d2";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"03a8") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"01ac";
        Y <= x"ab87";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"5625") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"2009";
        Y <= x"e814";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2008") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"2a24";
        Y <= x"2de1";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2de2") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"b438";
        Y <= x"efac";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"159c";
        Y <= x"5539";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ea64") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"79c1";
        Y <= x"9ba8";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"de19") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"8db2";
        Y <= x"e8ef";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"8db3") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"831a";
        Y <= x"1c98";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"d5b7";
        Y <= x"6f45";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"d8e7";
        Y <= x"9836";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"bf4f") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"4dc8";
        Y <= x"b887";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4779") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"9b92";
        Y <= x"2e4e";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"9b93") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"2cc2";
        Y <= x"27bb";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"547d") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"4275";
        Y <= x"b876";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"cf4d";
        Y <= x"6ef7";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"6ef8") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"dc9d";
        Y <= x"569c";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a963") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"7629";
        Y <= x"6eab";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"6eab") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"3d1f";
        Y <= x"9bd8";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"1005";
        Y <= x"48c7";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b738") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"d04c";
        Y <= x"991a";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"66e5") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"465c";
        Y <= x"aba5";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"aba4") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"3409";
        Y <= x"1d67";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"3408") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"5b5c";
        Y <= x"147d";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b921") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"75af";
        Y <= x"9d4b";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"75ae") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"61a6";
        Y <= x"d140";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"9066") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"8782";
        Y <= x"3f8f";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"406a";
        Y <= x"8054";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4069") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"df3f";
        Y <= x"b51c";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"df3e") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"6a86";
        Y <= x"0006";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"6a87") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"4fa5";
        Y <= x"cf09";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7f64") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"40be";
        Y <= x"7b88";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3aca") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"4290";
        Y <= x"0037";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4259") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"be71";
        Y <= x"fe89";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"fef9") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"8ddd";
        Y <= x"e670";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"bd24";
        Y <= x"5f16";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a0ea") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '1') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"e30b";
        Y <= x"603a";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"9fc5") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"7008";
        Y <= x"c38f";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"4ccb";
        Y <= x"890b";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b335") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"3c1b";
        Y <= x"b9f0";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"2328";
        Y <= x"9b04";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"dcd7") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"fed1";
        Y <= x"8889";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"89b8") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"768f";
        Y <= x"d8b4";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"febf") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"380e";
        Y <= x"3b8a";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"3b89") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"6292";
        Y <= x"31d2";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"6291") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"f862";
        Y <= x"7399";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"fbfb") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"f005";
        Y <= x"606c";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"8f99") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"f44c";
        Y <= x"246c";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"cfe0") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"ee48";
        Y <= x"0a88";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ee47") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"cd67";
        Y <= x"789b";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"cd68") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"5196";
        Y <= x"7ded";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"7ded") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"1df6";
        Y <= x"02d9";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"02d9") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"9c79";
        Y <= x"ee8b";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"8c09") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"2fb2";
        Y <= x"6ad6";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"d04d") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"dc4c";
        Y <= x"2158";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2158") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"4e85";
        Y <= x"1004";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"9b2a";
        Y <= x"415b";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"a798";
        Y <= x"f09e";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"a798") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"93c8";
        Y <= x"41fe";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ae36") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"b079";
        Y <= x"de34";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"8ead") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"52bd";
        Y <= x"6536";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4034") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"6498";
        Y <= x"38cc";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"38cd") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"f594";
        Y <= x"be14";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"c047";
        Y <= x"12af";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3fb8") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"e7d5";
        Y <= x"b729";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"182b") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"9667";
        Y <= x"acec";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"aceb") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"7619";
        Y <= x"1145";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"1001") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"7c1b";
        Y <= x"38c3";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"bca8") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"25cb";
        Y <= x"6ab0";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"da34") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"e261";
        Y <= x"9647";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e262") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"8970";
        Y <= x"3edd";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"8970") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"fc73";
        Y <= x"7dc9";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"8236") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"4ad5";
        Y <= x"a5b6";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f08b") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"85bb";
        Y <= x"2d99";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"85bb") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"b89a";
        Y <= x"f452";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3bb8") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"2d6a";
        Y <= x"3c80";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"ef9a";
        Y <= x"6d87";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ef99") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"49f3";
        Y <= x"ccdf";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"49f3") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"883d";
        Y <= x"ae1f";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ae3f") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"7613";
        Y <= x"ecd5";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7614") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"9e10";
        Y <= x"ffd0";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"9e11") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"ff0a";
        Y <= x"0826";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"00f5") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"30cc";
        Y <= x"c03f";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"c03e") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"8a47";
        Y <= x"1193";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"8a46") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"fd71";
        Y <= x"16f3";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"b927";
        Y <= x"5322";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"57cb";
        Y <= x"c85d";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"37a2") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"ea23";
        Y <= x"885d";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"885e") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"086c";
        Y <= x"4409";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4409") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"81bf";
        Y <= x"5ae4";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"6e19";
        Y <= x"d9b8";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2647") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"7410";
        Y <= x"2328";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2000") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"7190";
        Y <= x"aed1";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"718f") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"de8c";
        Y <= x"53ad";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"dfad") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"e992";
        Y <= x"2e08";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"e992") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"86b2";
        Y <= x"7992";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"272c";
        Y <= x"1477";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"2072";
        Y <= x"6daf";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4d3d") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"3734";
        Y <= x"ed07";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"c8cc") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"9def";
        Y <= x"c38a";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"da65") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"02b0";
        Y <= x"45f7";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"02af") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"db09";
        Y <= x"6687";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4201") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"2875";
        Y <= x"b71d";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2876") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"080f";
        Y <= x"7144";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"080e") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"6aaf";
        Y <= x"9c94";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"9551") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"4053";
        Y <= x"8dbf";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4054") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"4f84";
        Y <= x"7e36";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4f84") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"9717";
        Y <= x"a4bb";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f25c") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"8152";
        Y <= x"54db";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7ead") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"38cf";
        Y <= x"4fc5";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e90a") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"e8b7";
        Y <= x"43ca";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4082") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"deda";
        Y <= x"fa1d";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"05e2") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"af7c";
        Y <= x"7e11";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"7e10") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"0a27";
        Y <= x"d008";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"fe3a";
        Y <= x"4a66";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4a22") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"67f6";
        Y <= x"861b";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"980a") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"cd1a";
        Y <= x"6626";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ef3e") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"33af";
        Y <= x"6d74";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2124") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"9d0b";
        Y <= x"9889";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"a3d5";
        Y <= x"2dcf";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2dd0") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"ee2a";
        Y <= x"053e";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"f223";
        Y <= x"00d2";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ff2d") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"54b8";
        Y <= x"73d7";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"73d8") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"9e38";
        Y <= x"aa37";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f401") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"5838";
        Y <= x"7cf9";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7cfa") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"f339";
        Y <= x"1b0e";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"1b0e") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"93fa";
        Y <= x"b689";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4976") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"f2a3";
        Y <= x"87d4";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"782b") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"da15";
        Y <= x"3544";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"da14") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"a3ad";
        Y <= x"cd6b";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"a3ac") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"fa3b";
        Y <= x"b036";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b5fb") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"f6d4";
        Y <= x"4714";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b8ec") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '1') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"9817";
        Y <= x"17dd";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e822") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"61c7";
        Y <= x"da15";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"afa0";
        Y <= x"b94f";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"afa0") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"1ded";
        Y <= x"4564";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ba9c") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '1') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"6218";
        Y <= x"4ef4";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4ef4") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"5fa9";
        Y <= x"44aa";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a056") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"788d";
        Y <= x"2778";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2008") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"9cde";
        Y <= x"3904";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"6322") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"c7cb";
        Y <= x"e1ae";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e7ef") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"5e99";
        Y <= x"76d4";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"5e9a") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"4a72";
        Y <= x"a1a5";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ebf7") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"4921";
        Y <= x"5f06";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4920") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"d06c";
        Y <= x"cbde";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"c04c") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"9e4b";
        Y <= x"d90a";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"61b4") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"481d";
        Y <= x"70de";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"70dd") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"3454";
        Y <= x"0057";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"cbac") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"1c2b";
        Y <= x"1485";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"1c2b") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"ed5d";
        Y <= x"a91a";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"bbbd") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"2017";
        Y <= x"a931";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"56ce") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"6314";
        Y <= x"d26b";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"9ceb") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"aa53";
        Y <= x"1413";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"aa52") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"388c";
        Y <= x"0f97";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"388c") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"d81a";
        Y <= x"f9a3";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f9a2") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"bf66";
        Y <= x"61b6";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"5329";
        Y <= x"2be5";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"acd6") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"569b";
        Y <= x"04a8";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"56bb") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '0') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"1c80";
        Y <= x"0c41";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"efc1") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"2bd3";
        Y <= x"096f";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2bff") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '0') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"ed42";
        Y <= x"069b";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"069c") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"018e";
        Y <= x"8304";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"fe72") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"d903";
        Y <= x"1e89";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4586") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"c213";
        Y <= x"7923";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"7923") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"1f2f";
        Y <= x"b0f8";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"b0f7") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"e5b9";
        Y <= x"7a3f";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"6431";
        Y <= x"6566";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"6567") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"3d74";
        Y <= x"e429";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"e429") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"5bac";
        Y <= x"0c09";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"fc93";
        Y <= x"0bf6";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f409") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"c8d4";
        Y <= x"4038";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"090c") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"d513";
        Y <= x"eeb4";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"114b") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"5569";
        Y <= x"c4f8";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"7270";
        Y <= x"2a9d";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7afd") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '0') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"7fd3";
        Y <= x"e6ed";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"66c1") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"becf";
        Y <= x"f543";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"c98c") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"94c6";
        Y <= x"d940";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"bb86") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"9902";
        Y <= x"7d4b";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"66fd") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"85fe";
        Y <= x"8f23";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"85ff") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"ceef";
        Y <= x"7d3f";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"7d6b";
        Y <= x"e81f";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e820") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"9a8a";
        Y <= x"dd76";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2289") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"dec6";
        Y <= x"b205";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"8f5e";
        Y <= x"0a6f";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f590") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"1d82";
        Y <= x"6411";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"6411") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"fe8f";
        Y <= x"ce0a";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"cf7b") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"dfeb";
        Y <= x"d9a4";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2014") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"8369";
        Y <= x"13a9";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"93e9") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"3562";
        Y <= x"121a";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"3561") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"234c";
        Y <= x"d8ac";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b560") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"a011";
        Y <= x"baf1";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"a011") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"9f06";
        Y <= x"dd5a";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"60f9") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"0072";
        Y <= x"52c2";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"4458";
        Y <= x"e61a";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"1f6b";
        Y <= x"5ff2";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e094") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"1bec";
        Y <= x"00b1";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"00b0") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"75e8";
        Y <= x"71da";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"75e8") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"4ab3";
        Y <= x"1cc0";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"d298";
        Y <= x"2630";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2d68") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"6817";
        Y <= x"c1a7";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"29be") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"1136";
        Y <= x"10bb";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"21f1") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"594a";
        Y <= x"943c";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"5949") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"aa59";
        Y <= x"164c";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"be5d") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"9321";
        Y <= x"9205";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"fee4") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"4d3e";
        Y <= x"8708";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b2c2") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"9a24";
        Y <= x"f232";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"8c56") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"30ef";
        Y <= x"96ed";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"10ed") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"8e36";
        Y <= x"711b";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"8e36") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"4bbd";
        Y <= x"37e0";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"37e1") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"41c1";
        Y <= x"970e";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"41c2") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"874a";
        Y <= x"ca17";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"7c03";
        Y <= x"f4fb";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"7c02") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"1bc7";
        Y <= x"17b4";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"5c86";
        Y <= x"1815";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"1815") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"8018";
        Y <= x"3af5";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"bb0d") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"1d2a";
        Y <= x"e93a";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e93b") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"24b5";
        Y <= x"7971";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"db4b") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"1857";
        Y <= x"2c80";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e7a8") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"2e46";
        Y <= x"66ea";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"d1b9") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"7403";
        Y <= x"c491";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"3894") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"4cb0";
        Y <= x"e310";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4cb1") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"0f82";
        Y <= x"5806";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0802") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"e3f3";
        Y <= x"e8b6";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"e86b";
        Y <= x"6f01";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"8696") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"aa23";
        Y <= x"63c8";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"63c9") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"d2e3";
        Y <= x"e1be";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2d1d") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"5521";
        Y <= x"5386";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"0da0";
        Y <= x"9367";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0da0") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"644c";
        Y <= x"661a";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"644d") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"ba0f";
        Y <= x"2820";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2800") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"9f03";
        Y <= x"47de";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"5725") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"2f97";
        Y <= x"e334";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2f98") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"2e18";
        Y <= x"cd47";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"cd48") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"dfc7";
        Y <= x"5ae7";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"dfc7") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"f415";
        Y <= x"5c5f";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f414") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"6ca9";
        Y <= x"3126";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"6ca8") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"5975";
        Y <= x"a2ec";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"1ae8";
        Y <= x"dde6";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"1ae9") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"adae";
        Y <= x"84c4";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"84c3") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '1') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"ebcb";
        Y <= x"71aa";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"1434") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"ef7a";
        Y <= x"4756";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4752") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"cbb0";
        Y <= x"e01c";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"abcc") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"dc55";
        Y <= x"535d";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2fb2") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"52b4";
        Y <= x"116b";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"f47f";
        Y <= x"3ee2";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f47e") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"c567";
        Y <= x"5aac";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"dfef") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"4da8";
        Y <= x"f4c1";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"0b84";
        Y <= x"8a6e";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"8a6f") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"1fb2";
        Y <= x"5b6f";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"1fb2") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"7f13";
        Y <= x"d6e2";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"57cf") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"de9a";
        Y <= x"94e9";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"af81";
        Y <= x"43e9";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"90fc";
        Y <= x"b68b";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"6f03") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"4b33";
        Y <= x"4769";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b896") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"b3f0";
        Y <= x"d1d6";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b3f1") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"91ac";
        Y <= x"323a";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"323a") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"f514";
        Y <= x"be08";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ff1c") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"b9b6";
        Y <= x"2072";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"df8d") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"68d6";
        Y <= x"7b56";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7bd6") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '0') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"0d13";
        Y <= x"8c9f";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0d12") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"306f";
        Y <= x"6956";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"99c5") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"8050";
        Y <= x"738c";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"738d") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"596c";
        Y <= x"9e9a";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"6166") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"4ff5";
        Y <= x"8c15";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4ff4") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"a3bd";
        Y <= x"3294";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"54cc";
        Y <= x"c0ca";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"54cc") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"c092";
        Y <= x"4989";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7709") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"c470";
        Y <= x"9070";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"be2a";
        Y <= x"c892";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"ae73";
        Y <= x"1599";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0411") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"0943";
        Y <= x"3714";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f6bc") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"23cc";
        Y <= x"14c4";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"dc33") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"313f";
        Y <= x"3b46";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"3106") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"40e3";
        Y <= x"4cc3";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b33c") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"c210";
        Y <= x"a33a";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"8d88";
        Y <= x"631f";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"e450";
        Y <= x"0d01";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"31c2";
        Y <= x"d459";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ce3e") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"9bc8";
        Y <= x"950a";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"06be") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"e229";
        Y <= x"098e";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0008") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"1dcc";
        Y <= x"ee36";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0c02") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"4735";
        Y <= x"15b5";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"d3cc";
        Y <= x"9253";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"3ebf";
        Y <= x"3c78";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3eff") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '0') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"2159";
        Y <= x"b8a0";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2000") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"4907";
        Y <= x"9822";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4f1b") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"b008";
        Y <= x"2839";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2838") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"dbd0";
        Y <= x"5f1d";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"dbcf") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"0b70";
        Y <= x"cb9d";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"922e";
        Y <= x"cf3d";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"822c") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"40e8";
        Y <= x"460c";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"804b";
        Y <= x"cdf0";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"3210") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '0') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"0f41";
        Y <= x"2007";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f0bf") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"1508";
        Y <= x"0c80";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"acf1";
        Y <= x"3820";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"530e") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '0') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"3567";
        Y <= x"10f2";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"1062") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"fe3d";
        Y <= x"da57";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"dc1a") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"a283";
        Y <= x"3705";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"a283") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '1') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"a606";
        Y <= x"74ac";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"74ab") report "Error in outcome (dec y)" severity note;
        assert (zr = '0') report "Error in zero flag (dec y)" severity note;
        assert (ng = '0') report "Error in negative flag (dec y)" severity note;
        wait for 1 ns;

        X <= x"4764";
        Y <= x"2cfa";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2cfa") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"bb86";
        Y <= x"05ae";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"bb85") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"1f60";
        Y <= x"635a";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"c973";
        Y <= x"ca0a";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"c972") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"78fb";
        Y <= x"dd76";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"dd76") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"f61f";
        Y <= x"825d";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"825e") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"cfab";
        Y <= x"ad60";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ddb5") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"c178";
        Y <= x"459d";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ba63") report "Error in outcome (minus y)" severity note;
        assert (zr = '0') report "Error in zero flag (minus y)" severity note;
        assert (ng = '1') report "Error in negative flag (minus y)" severity note;
        wait for 1 ns;

        X <= x"33f4";
        Y <= x"945d";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"33f5") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"077b";
        Y <= x"5643";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"4ec8") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"d007";
        Y <= x"4aef";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b510") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"5113";
        Y <= x"b034";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"1010") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"5680";
        Y <= x"b41a";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a266") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"8987";
        Y <= x"0a75";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7679") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"7307";
        Y <= x"92c0";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"92c1") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"bcd0";
        Y <= x"ad23";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"bdf3") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"510a";
        Y <= x"06ff";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"57ff") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '0') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"8902";
        Y <= x"6f59";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"e657") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"e573";
        Y <= x"ec41";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"b61b";
        Y <= x"e403";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"49e5") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"2762";
        Y <= x"f4e3";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"1c45") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"9752";
        Y <= x"61d1";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"865d";
        Y <= x"3360";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"3360") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '0') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"9076";
        Y <= x"4c6f";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"96ed";
        Y <= x"ca2c";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"822c") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"b077";
        Y <= x"3ab4";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"b076") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"a3c7";
        Y <= x"2f09";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"8b42") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"3314";
        Y <= x"52b7";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"52b8") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '0') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"bdd7";
        Y <= x"9c0f";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"de38") report "Error in outcome (sub_yx)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_yx)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_yx)" severity note;
        wait for 1 ns;

        X <= x"58aa";
        Y <= x"48d4";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"3a4b";
        Y <= x"c60a";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"7441") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '0') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"b34f";
        Y <= x"1350";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b350") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"a1fd";
        Y <= x"b16b";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b16c") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"5b2b";
        Y <= x"9ded";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"f918") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"ac38";
        Y <= x"1d22";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ac37") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '1') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"1a3d";
        Y <= x"6e1b";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"ac22") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"7e8e";
        Y <= x"3942";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"7e8e") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"0728";
        Y <= x"2723";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"c69b";
        Y <= x"152b";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"20c4";
        Y <= x"0b1e";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"2bde") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '0') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"a88f";
        Y <= x"7277";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"a890") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '1') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"8ae9";
        Y <= x"55e5";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"aa1a") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '1') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"6ff5";
        Y <= x"0e7d";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"ba65";
        Y <= x"742f";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"2e94") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"76a4";
        Y <= x"b36f";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"b36f") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"f9e3";
        Y <= x"4653";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"061d") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '0') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"82c6";
        Y <= x"5360";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"6137";
        Y <= x"a0b0";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"7976";
        Y <= x"8f9a";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"cac0";
        Y <= x"847b";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"cefb") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"9354";
        Y <= x"c3c2";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"8340") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"d22f";
        Y <= x"759e";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f7bf") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"3bcb";
        Y <= x"d697";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"d697") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"236d";
        Y <= x"31ad";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"551a") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '0') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"a97f";
        Y <= x"6349";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"eb7f") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"171a";
        Y <= x"d188";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"e8a2") report "Error in outcome (add)" severity note;
        assert (zr = '0') report "Error in zero flag (add)" severity note;
        assert (ng = '1') report "Error in negative flag (add)" severity note;
        wait for 1 ns;

        X <= x"9852";
        Y <= x"d426";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"c42c") report "Error in outcome (sub_xy)" severity note;
        assert (zr = '0') report "Error in zero flag (sub_xy)" severity note;
        assert (ng = '1') report "Error in negative flag (sub_xy)" severity note;
        wait for 1 ns;

        X <= x"6984";
        Y <= x"c523";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"967c") report "Error in outcome (minus x)" severity note;
        assert (zr = '0') report "Error in zero flag (minus x)" severity note;
        assert (ng = '1') report "Error in negative flag (minus x)" severity note;
        wait for 1 ns;

        X <= x"611b";
        Y <= x"4d43";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"611c") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"e662";
        Y <= x"54c5";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"d285";
        Y <= x"35e7";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;

        X <= x"9b95";
        Y <= x"eef0";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"eef0") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"37b8";
        Y <= x"9d51";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"62ae") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"d5b1";
        Y <= x"233b";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"5771";
        Y <= x"a3b3";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"5770") report "Error in outcome (dec x)" severity note;
        assert (zr = '0') report "Error in zero flag (dec x)" severity note;
        assert (ng = '0') report "Error in negative flag (dec x)" severity note;
        wait for 1 ns;

        X <= x"01a2";
        Y <= x"b969";
        zx <= '0';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"01a3") report "Error in outcome (inc x)" severity note;
        assert (zr = '0') report "Error in zero flag (inc x)" severity note;
        assert (ng = '0') report "Error in negative flag (inc x)" severity note;
        wait for 1 ns;

        X <= x"c45d";
        Y <= x"8d12";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"72ed") report "Error in outcome (not y)" severity note;
        assert (zr = '0') report "Error in zero flag (not y)" severity note;
        assert (ng = '0') report "Error in negative flag (not y)" severity note;
        wait for 1 ns;

        X <= x"1689";
        Y <= x"9959";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"1689") report "Error in outcome (x)" severity note;
        assert (zr = '0') report "Error in zero flag (x)" severity note;
        assert (ng = '0') report "Error in negative flag (x)" severity note;
        wait for 1 ns;

        X <= x"f471";
        Y <= x"63b4";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"4151";
        Y <= x"4219";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"4011") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '0') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"6d3d";
        Y <= x"2c02";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"dc74";
        Y <= x"86e8";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"86e9") report "Error in outcome (inc y)" severity note;
        assert (zr = '0') report "Error in zero flag (inc y)" severity note;
        assert (ng = '1') report "Error in negative flag (inc y)" severity note;
        wait for 1 ns;

        X <= x"9212";
        Y <= x"2d8b";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"6f11";
        Y <= x"db68";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"db68") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"cc8b";
        Y <= x"c345";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"c001") report "Error in outcome (and)" severity note;
        assert (zr = '0') report "Error in zero flag (and)" severity note;
        assert (ng = '1') report "Error in negative flag (and)" severity note;
        wait for 1 ns;

        X <= x"dd9d";
        Y <= x"b168";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"15fb";
        Y <= x"9b20";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"ffff") report "Error in outcome (minus one)" severity note;
        assert (zr = '0') report "Error in zero flag (minus one)" severity note;
        assert (ng = '1') report "Error in negative flag (minus one)" severity note;
        wait for 1 ns;

        X <= x"4b89";
        Y <= x"7a5b";
        zx <= '0';
        zy <= '1';
        nx <= '0';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"b476") report "Error in outcome (not x)" severity note;
        assert (zr = '0') report "Error in zero flag (not x)" severity note;
        assert (ng = '1') report "Error in negative flag(not x)" severity note;
        wait for 1 ns;

        X <= x"b6a0";
        Y <= x"1f7e";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"bffe") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"f0b2";
        Y <= x"a442";
        zx <= '1';
        zy <= '1';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"0000") report "Error in outcome (zero)" severity note;
        assert (zr = '1') report "Error in zero flag (zero)" severity note;
        assert (ng = '0') report "Error in negative flag (zero)" severity note;
        wait for 1 ns;

        X <= x"f5dc";
        Y <= x"f3fc";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"f7fc") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"4eeb";
        Y <= x"e4ba";
        zx <= '1';
        zy <= '0';
        nx <= '1';
        ny <= '0';
        f <= '0';
        no <= '0';
        wait for 1 ns;
        assert (Z = x"e4ba") report "Error in outcome (y)" severity note;
        assert (zr = '0') report "Error in zero flag (y)" severity note;
        assert (ng = '1') report "Error in negative flag (y)" severity note;
        wait for 1 ns;

        X <= x"d7b2";
        Y <= x"4e81";
        zx <= '0';
        zy <= '0';
        nx <= '1';
        ny <= '1';
        f <= '0';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"dfb3") report "Error in outcome (or)" severity note;
        assert (zr = '0') report "Error in zero flag (or)" severity note;
        assert (ng = '1') report "Error in negative flag (or)" severity note;
        wait for 1 ns;

        X <= x"91c9";
        Y <= x"80e6";
        zx <= '1';
        zy <= '1';
        nx <= '1';
        ny <= '1';
        f <= '1';
        no <= '1';
        wait for 1 ns;
        assert (Z = x"0001") report "Error in outcome (one)" severity note;
        assert (zr = '0') report "Error in zero flag (one)" severity note;
        assert (ng = '0') report "Error in negative flag (one)" severity note;
        wait for 1 ns;



        report "Simulation done";

        wait;
    end process;


    -------------------------------------------------------------------------------
    -- DUT
    -------------------------------------------------------------------------------
    DUT: component alu port map(
        X => X,
        Y => Y,
        Z => Z,
        zx => zx,
        zy => zy,
        nx => nx,
        ny => ny,
        f => f,
        no => no,
        zr => zr,
        ng => ng
    );

end Behavioural;
