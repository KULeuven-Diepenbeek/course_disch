    PSTIM: process
    begin
        X <= x"C";
        Y <= x"3";
        zx <= '0';
        zy <= '0';
        nx <= '0';
        ny <= '0';
        f <= '1';
        no <= '0';

        wait;
    end process;