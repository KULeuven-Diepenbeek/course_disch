library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity alu_tb is
end entity alu_tb;

architecture Behavioural of alu_tb is
    component alu is
        port(
            operand1 : in std_logic_vector(32-1 downto 0);
            operand2 : in std_logic_vector(32-1 downto 0);
            ALUOp : in std_logic_vector(2 downto 0);
            arith_logic_b : in STD_LOGIC;
            signed_unsigned_b : in STD_LOGIC;
            result : out std_logic_vector(32-1 downto 0);
            equal : out STD_LOGIC;
            x_lt_y_u : out STD_LOGIC;
            x_lt_y_s : out STD_LOGIC
        );
    end component alu;

    signal operand1 : std_logic_vector(32-1 downto 0);
    signal operand2 : std_logic_vector(32-1 downto 0);
    signal ALUOp : std_logic_vector(2 downto 0);
    signal arith_logic_b : STD_LOGIC;
    signal signed_unsigned_b : STD_LOGIC;
    signal result : std_logic_vector(32-1 downto 0);
    signal equal : STD_LOGIC;
    signal x_lt_y_u : STD_LOGIC;
    signal x_lt_y_s : STD_LOGIC;

begin

    PSTIM: process
        variable good_checks : natural;
        variable bad_checks : natural;
    begin
        operand1 <= (others => '0');
        operand2 <= (others => '0');
        ALUOp <= (others => '0');
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        good_checks := 0;
        bad_checks := 0;
        wait for 4 ns;

        -- apply stimuli
        operand1 <= x"8ffb9e07"; -- 2415631879
        operand2 <= x"fdcea5ee"; -- 4258178542
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8dca8406" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"88abdb82"; -- 2292964226
        operand2 <= x"0328f349"; -- 53015369
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0028d300" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f2c9d056"; -- 4073312342
        operand2 <= x"27205659"; -- 656430681
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"22005050" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ca6eed1b"; -- 3396267291
        operand2 <= x"226a7a5a"; -- 577403482
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"026a681a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"31a45d63"; -- 832855395
        operand2 <= x"9ede3f43"; -- 2665365315
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"10841d43" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9ff5826b"; -- 2683667051
        operand2 <= x"3dd4f32a"; -- 1037366058
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1dd4822a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3a84fa2a"; -- 981793322
        operand2 <= x"15391e3d"; -- 356064829
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"10001a28" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"eede221f"; -- 4007535135
        operand2 <= x"2c832a54"; -- 746793556
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2c822214" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"703ae0cb"; -- 1882906827
        operand2 <= x"4e1ce0dd"; -- 1310515421
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4018e0c9" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"07f588d6"; -- 133531862
        operand2 <= x"f30be11b"; -- 4077642011
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"03018012" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"16405e10"; -- 373317136
        operand2 <= x"64c1129a"; -- 1690374810
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"04401210" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2744478f"; -- 658786191
        operand2 <= x"f709e610"; -- 4144621072
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"27004600" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"62288a24"; -- 1646823972
        operand2 <= x"7c8968cd"; -- 2089380045
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"60080804" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b6d13a3d"; -- 3067165245
        operand2 <= x"3039489f"; -- 809060511
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3011081d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"93004497"; -- 2466268311
        operand2 <= x"5e96822f"; -- 1586922031
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"12000007" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"64cd1da1"; -- 1691164065
        operand2 <= x"624cac2a"; -- 1649191978
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"604c0c20" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"64accc7b"; -- 1689046139
        operand2 <= x"f5349651"; -- 4113864273
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"64248451" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b12118dd"; -- 2971736285
        operand2 <= x"92723b16"; -- 2456959766
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"90201814" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0b54582f"; -- 190076975
        operand2 <= x"32846f92"; -- 847540114
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"02044802" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1959fdff"; -- 425328127
        operand2 <= x"b7a97080"; -- 3081334912
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"11097080" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4687005f"; -- 1183252575
        operand2 <= x"de7568dd"; -- 3732236509
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4605005d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7ce8d0b7"; -- 2095632567
        operand2 <= x"9c37405e"; -- 2620866654
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1c204016" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1e6e1816"; -- 510531606
        operand2 <= x"4bbfa955"; -- 1270851925
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0a2e0814" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1a60fff2"; -- 442564594
        operand2 <= x"47fd8e38"; -- 1207799352
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"02608e30" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bc469dcb"; -- 3158744523
        operand2 <= x"ae2b2726"; -- 2922063654
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ac020502" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"22220917"; -- 572655895
        operand2 <= x"3113dcae"; -- 823385262
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"20020806" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dc3ab18a"; -- 3694834058
        operand2 <= x"e7f11049"; -- 3891335241
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c4301008" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5ccb26a8"; -- 1556817576
        operand2 <= x"e37deb1c"; -- 3816680220
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"40492208" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"16f82f82"; -- 385363842
        operand2 <= x"2d3ffbf4"; -- 759167988
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"04382b80" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8f40b5ad"; -- 2403382701
        operand2 <= x"ac67ab12"; -- 2892475154
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8c40a100" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2a9cab40"; -- 714910528
        operand2 <= x"b279b9f0"; -- 2994321904
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2218a940" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"54c2722b"; -- 1422029355
        operand2 <= x"12239cac"; -- 304323756
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"10021028" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"475cb186"; -- 1197257094
        operand2 <= x"56c34fac"; -- 1455640492
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"46400184" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b163c7c7"; -- 2976106439
        operand2 <= x"b79cbe57"; -- 3080502871
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b1008647" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"65ec779d"; -- 1709995933
        operand2 <= x"00750cc0"; -- 7670976
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00640480" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"57382652"; -- 1463297618
        operand2 <= x"798958d3"; -- 2039044307
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"51080052" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6e3062b8"; -- 1848664760
        operand2 <= x"78619c12"; -- 2019662866
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"68200010" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c829c53a"; -- 3358180666
        operand2 <= x"beff4ed8"; -- 3204402904
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"88294418" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f3bb0de3"; -- 4089122275
        operand2 <= x"85dd59bc"; -- 2245876156
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"819909a0" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a5147e16"; -- 2769583638
        operand2 <= x"1797bc1c"; -- 395820060
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"05143c14" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b3e57c71"; -- 3018161265
        operand2 <= x"8fbe14c4"; -- 2411599044
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"83a41440" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"42c150f2"; -- 1119965426
        operand2 <= x"fcb0ec42"; -- 4239453250
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"40804042" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2535bb06"; -- 624278278
        operand2 <= x"aa072ce9"; -- 2852596969
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"20052800" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"58a69364"; -- 1487311716
        operand2 <= x"c3a4743c"; -- 3282334780
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"40a41024" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"503fc5fc"; -- 1346356732
        operand2 <= x"dfe511cd"; -- 3756331469
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"502501cc" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"76ad514a"; -- 1991070026
        operand2 <= x"d1288753"; -- 3509094227
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"50280142" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"83c827d9"; -- 2210932697
        operand2 <= x"0088be43"; -- 8961603
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00882641" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e6788de3"; -- 3866660323
        operand2 <= x"5f813599"; -- 1602303385
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"46000581" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4965d65b"; -- 1231410779
        operand2 <= x"60aea946"; -- 1622059334
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"40248042" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5e211b6e"; -- 1579228014
        operand2 <= x"c12f262d"; -- 3241092653
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4021022c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"20e7676b"; -- 552036203
        operand2 <= x"4ff0176b"; -- 1341134699
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00e0076b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f6a98b7d"; -- 4138306429
        operand2 <= x"27f8f66c"; -- 670627436
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"26a8826c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5dce5345"; -- 1573802821
        operand2 <= x"8583f403"; -- 2240017411
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"05825001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a4dee0eb"; -- 2766069995
        operand2 <= x"634941ef"; -- 1665745391
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"204840eb" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"53dc88b4"; -- 1406961844
        operand2 <= x"c5b4c863"; -- 3316959331
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"41948820" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d436e8f1"; -- 3560368369
        operand2 <= x"6b0da91b"; -- 1796057371
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4004a811" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5ef16aff"; -- 1592879871
        operand2 <= x"5dc5256c"; -- 1573201260
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"5cc1206c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8b1420c2"; -- 2333352130
        operand2 <= x"ba8fec3f"; -- 3129994303
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8a042002" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"23bbd941"; -- 599513409
        operand2 <= x"63267d94"; -- 1663466900
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"23225900" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5f4cdc6a"; -- 1598872682
        operand2 <= x"a8a9365e"; -- 2829661790
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0808144a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6a427569"; -- 1782740329
        operand2 <= x"892cf5a4"; -- 2301425060
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"08007520" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d204761d"; -- 3523507741
        operand2 <= x"4328408a"; -- 1126711434
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"42004008" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8beb61c2"; -- 2347459010
        operand2 <= x"eddd8cce"; -- 3990719694
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"89c900c2" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"218f9bc6"; -- 563059654
        operand2 <= x"54e3f7d4"; -- 1424226260
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"008393c4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dd05498b"; -- 3708111243
        operand2 <= x"df299d42"; -- 3744046402
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"dd010902" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dfaa3312"; -- 3752473362
        operand2 <= x"76af7e86"; -- 1991212678
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"56aa3202" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"da9a2f9c"; -- 3667537820
        operand2 <= x"870e1e31"; -- 2265849393
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"820a0e10" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e1db5efe"; -- 3789250302
        operand2 <= x"344546f8"; -- 876955384
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"204146f8" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"144ce8e8"; -- 340584680
        operand2 <= x"e078784a"; -- 3765991498
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00486848" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4c514ce6"; -- 1280396518
        operand2 <= x"9492984b"; -- 2492635211
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"04100842" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5d879191"; -- 1569165713
        operand2 <= x"c3bb3e25"; -- 3283828261
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"41831001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e0f755ea"; -- 3774305770
        operand2 <= x"cbf5071f"; -- 3421832991
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c0f5050a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d31c0fad"; -- 3541831597
        operand2 <= x"654b613d"; -- 1699438909
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4108012d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8c5156b2"; -- 2354140850
        operand2 <= x"630d2f64"; -- 1661808484
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00010620" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"481ea14d"; -- 1209966925
        operand2 <= x"97290bf8"; -- 2536049656
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00080148" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b267cbb7"; -- 2993146807
        operand2 <= x"835d467e"; -- 2203928190
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"82454236" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"239fe57d"; -- 597681533
        operand2 <= x"58ffb849"; -- 1493153865
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"009fa049" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"58b026fb"; -- 1487939323
        operand2 <= x"d0a4046e"; -- 3500409966
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"50a0046a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8cd5e783"; -- 2362828675
        operand2 <= x"7a48078b"; -- 2051540875
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"08400783" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"07db6fd1"; -- 131821521
        operand2 <= x"d5a97e39"; -- 3584654905
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"05896e11" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8c7771cb"; -- 2356638155
        operand2 <= x"e7f3044b"; -- 3891463243
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8473004b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7f1ecefd"; -- 2132725501
        operand2 <= x"c9a7b4d3"; -- 3383211219
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"490684d1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"05cbf29c"; -- 97251996
        operand2 <= x"0aad1c36"; -- 179117110
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00891014" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"66e70a98"; -- 1726417560
        operand2 <= x"381c189b"; -- 941365403
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"20040898" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"34efd566"; -- 888132966
        operand2 <= x"7a26f016"; -- 2049372182
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3026d006" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d9cd13ea"; -- 3654095850
        operand2 <= x"6fbdd037"; -- 1874710583
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"498d1022" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4cf4834d"; -- 1291092813
        operand2 <= x"e7e8407d"; -- 3890757757
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"44e0004d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c7f71e77"; -- 3354861175
        operand2 <= x"203ff97e"; -- 541063550
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00371876" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c61a1b78"; -- 3323599736
        operand2 <= x"aa6257e8"; -- 2858571752
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"82021368" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"115cea8a"; -- 291302026
        operand2 <= x"4efd2da1"; -- 1325215137
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"005c2880" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9d6eed29"; -- 2641292585
        operand2 <= x"f6a3f89c"; -- 4137941148
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9422e808" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"99aee5d3"; -- 2578376147
        operand2 <= x"def41859"; -- 3740538969
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"98a40051" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9387d355"; -- 2475152213
        operand2 <= x"a10257d2"; -- 2701285330
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"81025350" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ea82e612"; -- 3934447122
        operand2 <= x"a5200b20"; -- 2770340640
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a0000200" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ec430721"; -- 3963815713
        operand2 <= x"d26deaef"; -- 3530418927
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c0410221" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"62fe6d94"; -- 1660841364
        operand2 <= x"c73f71d1"; -- 3342823889
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"423e6190" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"cfa9f920"; -- 3484023072
        operand2 <= x"b598c383"; -- 3046687619
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8588c100" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"57ce2cde"; -- 1473129694
        operand2 <= x"37df90aa"; -- 937398442
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"17ce008a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0bb4d7b9"; -- 196401081
        operand2 <= x"a02ea5b9"; -- 2687411641
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"002485b9" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"327a4a09"; -- 846875145
        operand2 <= x"04fd76f0"; -- 83719920
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00784200" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"28f6b2e9"; -- 687256297
        operand2 <= x"43404b16"; -- 1128286998
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00400200" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b1fa43c6"; -- 2985968582
        operand2 <= x"1000b087"; -- 268480647
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"10000086" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8a9c6526"; -- 2325505318
        operand2 <= x"05c9ae9a"; -- 97103514
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00882402" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6f7284e0"; -- 1869776096
        operand2 <= x"385edd65"; -- 945741157
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"28528460" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c06fb5f8"; -- 3228546552
        operand2 <= x"10a975fe"; -- 279541246
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"002935f8" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"997a718b"; -- 2574938507
        operand2 <= x"3fc5c8ea"; -- 1069926634
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1940408a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4a1d828e"; -- 1243447950
        operand2 <= x"49617e8f"; -- 1231126159
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4801028e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"89cbb370"; -- 2311828336
        operand2 <= x"1e2389cc"; -- 505645516
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"08038140" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fabd687c"; -- 4206717052
        operand2 <= x"695af366"; -- 1767568230
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"68186064" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"23d6c9fd"; -- 601278973
        operand2 <= x"2868c9d4"; -- 677956052
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2040c9d4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"48f76749"; -- 1224173385
        operand2 <= x"18dcaaf1"; -- 417114865
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"08d42241" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"297c7c34"; -- 696024116
        operand2 <= x"67d72d5d"; -- 1742155101
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"21542c14" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d69dcf5a"; -- 3600666458
        operand2 <= x"e142ece9"; -- 3779259625
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c000cc48" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"374f0d63"; -- 927927651
        operand2 <= x"7a0d6a3d"; -- 2047699517
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"320d0821" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"835968ba"; -- 2203674810
        operand2 <= x"1c56920d"; -- 475435533
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00500008" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e94a5e2d"; -- 3913965101
        operand2 <= x"8bcea9af"; -- 2345576879
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"894a082d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d41f3e9f"; -- 3558817439
        operand2 <= x"3cc0951f"; -- 1019254047
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1400141f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"058d2024"; -- 93134884
        operand2 <= x"ba8d78ef"; -- 3129833711
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"008d2024" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0d58775c"; -- 223901532
        operand2 <= x"f6a09ffc"; -- 4137721852
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0400175c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"017c5c48"; -- 24927304
        operand2 <= x"825a7cec"; -- 2186968300
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00585c48" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"189100cd"; -- 412156109
        operand2 <= x"fdc7d53b"; -- 4257731899
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"18810009" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d0d2d1c7"; -- 3503477191
        operand2 <= x"f6e249e6"; -- 4142025190
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d0c241c6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"21140678"; -- 554960504
        operand2 <= x"3cba5e1d"; -- 1018846749
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"20100618" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c092f8d8"; -- 3230857432
        operand2 <= x"de88a52a"; -- 3733497130
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c080a008" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9775d938"; -- 2541082936
        operand2 <= x"f4b58517"; -- 4105536791
        ALUOp <= "000";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"94358110" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"13d23990"; -- 332544400
        operand2 <= x"47936732"; -- 1200842546
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"57d37fb2" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f93f1373"; -- 4181660531
        operand2 <= x"c13675a6"; -- 3241571750
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f93f77f7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5d9c3bff"; -- 1570520063
        operand2 <= x"b69aad81"; -- 3063590273
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ff9ebfff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e1173cd6"; -- 3776396502
        operand2 <= x"1bc1aab6"; -- 465676982
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fbd7bef6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"463a2a42"; -- 1178217026
        operand2 <= x"e0338126"; -- 3761471782
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"e63bab66" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"188af80a"; -- 411760650
        operand2 <= x"dec8ca1d"; -- 3737700893
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"decafa1f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fabe8138"; -- 4206788920
        operand2 <= x"57c31b8f"; -- 1472404367
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffff9bbf" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c57e4ecd"; -- 3313389261
        operand2 <= x"ecc24b01"; -- 3972156161
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"edfe4fcd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e739a2a3"; -- 3879314083
        operand2 <= x"f8f0ffce"; -- 4176543694
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fff9ffef" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"29e28bcd"; -- 702712781
        operand2 <= x"f768c8c4"; -- 4150839492
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffeacbcd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d72bc906"; -- 3609970950
        operand2 <= x"1abc488d"; -- 448546957
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"dfbfc98f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e417e295"; -- 3826770581
        operand2 <= x"7fe0a75e"; -- 2145429342
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fff7e7df" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"039a8788"; -- 60458888
        operand2 <= x"b67da85e"; -- 3061688414
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b7ffafde" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5c38a64b"; -- 1547216459
        operand2 <= x"2d9dc3ae"; -- 765313966
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7dbde7ef" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d526892a"; -- 3576072490
        operand2 <= x"04c6b4a5"; -- 80131237
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d5e6bdaf" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"47ab5904"; -- 1202411780
        operand2 <= x"2f764ea2"; -- 796282530
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6fff5fa6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e0729687"; -- 3765606023
        operand2 <= x"389e1954"; -- 949885268
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f8fe9fd7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"11dbd77d"; -- 299620221
        operand2 <= x"b30526dc"; -- 3003459292
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b3dff7fd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"34106c42"; -- 873491522
        operand2 <= x"60f82bb2"; -- 1626876850
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"74f86ff2" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e680255d"; -- 3867157853
        operand2 <= x"48a67f96"; -- 1218871190
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"eea67fdf" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"eec12b9f"; -- 4005637023
        operand2 <= x"57add324"; -- 1471009572
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffedfbbf" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"572a163e"; -- 1462375998
        operand2 <= x"f8837278"; -- 4169364088
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffab767e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b7b745d2"; -- 3082241490
        operand2 <= x"e76e0b29"; -- 3882748713
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f7ff4ffb" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dceade68"; -- 3706379880
        operand2 <= x"fc57a1f2"; -- 4233601522
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fcfffffa" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ba1a22eb"; -- 3122275051
        operand2 <= x"e69eebd6"; -- 3869174742
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fe9eebff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ccb65d42"; -- 3434503490
        operand2 <= x"c424bfcc"; -- 3290742732
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ccb6ffce" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1c5f617a"; -- 476012922
        operand2 <= x"a14386fe"; -- 2705557246
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bd5fe7fe" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"88538444"; -- 2287174724
        operand2 <= x"bbf8cad1"; -- 3153644241
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bbfbced5" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8414cbf2"; -- 2215955442
        operand2 <= x"15fa78cd"; -- 368736461
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"95fefbff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7a0eb403"; -- 2047783939
        operand2 <= x"a66a9413"; -- 2792002579
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fe6eb413" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3f7e1361"; -- 1065227105
        operand2 <= x"0915d30c"; -- 152425228
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3f7fd36d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2240202a"; -- 574627882
        operand2 <= x"dc20ffff"; -- 3693150207
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fe60ffff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"620b3623"; -- 1644901923
        operand2 <= x"3dc189b9"; -- 1036093881
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7fcbbfbb" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"26c37b6f"; -- 650345327
        operand2 <= x"8d69c089"; -- 2372518025
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"afebfbef" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1d000d93"; -- 486542739
        operand2 <= x"24fcf883"; -- 620558467
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3dfcfd93" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bbe264eb"; -- 3152176363
        operand2 <= x"806c2c70"; -- 2154572912
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bbee6cfb" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"46f42d4a"; -- 1190407498
        operand2 <= x"0a3d1014"; -- 171773972
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4efd3d5e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a2055286"; -- 2718257798
        operand2 <= x"dbb0d787"; -- 3685799815
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fbb5d787" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d6657ce3"; -- 3596975331
        operand2 <= x"8e2373ef"; -- 2384688111
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"de677fef" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9ec639bb"; -- 2663791035
        operand2 <= x"22a94dba"; -- 581520826
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"beef7dbb" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"43378657"; -- 1127712343
        operand2 <= x"60a6b642"; -- 1621538370
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"63b7b657" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9f7040c3"; -- 2674933955
        operand2 <= x"8faece44"; -- 2410597956
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9ffecec7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"180c8200"; -- 403472896
        operand2 <= x"abfa5590"; -- 2885309840
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bbfed790" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f5cdf443"; -- 4123915331
        operand2 <= x"1e8e49be"; -- 512641470
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffcffdff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"055ea2db"; -- 90088155
        operand2 <= x"7d545cbb"; -- 2102680763
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7d5efefb" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6b388a25"; -- 1798867493
        operand2 <= x"8f52a43f"; -- 2404557887
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ef7aae3f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3adde279"; -- 987619961
        operand2 <= x"3eb84096"; -- 1052262550
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3efde2ff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"39481b53"; -- 961026899
        operand2 <= x"5b0ef0b1"; -- 1527705777
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7b4efbf3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4bcf6236"; -- 1271882294
        operand2 <= x"96102aea"; -- 2517641962
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"dfdf6afe" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"003f95b3"; -- 4167091
        operand2 <= x"2bf8e06d"; -- 737730669
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2bfff5ff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7e8954a5"; -- 2122929317
        operand2 <= x"5325e6c8"; -- 1394992840
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7fadf6ed" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8039de9b"; -- 2151276187
        operand2 <= x"aa768f6f"; -- 2859896687
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"aa7fdfff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0e0ded9d"; -- 235793821
        operand2 <= x"b57af5e4"; -- 3044734436
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bf7ffdfd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"90f23aa5"; -- 2431793829
        operand2 <= x"29c73733"; -- 700921651
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b9f73fb7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e04003fd"; -- 3762291709
        operand2 <= x"773c9523"; -- 2000459043
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f77c97ff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d612e98f"; -- 3591563663
        operand2 <= x"438d6eae"; -- 1133342382
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d79fefaf" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3ece04cd"; -- 1053689037
        operand2 <= x"529d0922"; -- 1386023202
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7edf0def" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"df821720"; -- 3749844768
        operand2 <= x"85bdf0eb"; -- 2243817707
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"dfbff7eb" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3ec811e4"; -- 1053299172
        operand2 <= x"3ffd9c07"; -- 1073585159
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3ffd9de7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"64ef76ac"; -- 1693415084
        operand2 <= x"d583ec5e"; -- 3582192734
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f5effefe" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"60d8456f"; -- 1624786287
        operand2 <= x"a04de360"; -- 2689459040
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"e0dde76f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"12828a13"; -- 310544915
        operand2 <= x"3ed78aa8"; -- 1054313128
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3ed78abb" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"37f5a8c1"; -- 938846401
        operand2 <= x"aefc4f03"; -- 2935770883
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bffdefc3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5317cc04"; -- 1394068484
        operand2 <= x"ac025820"; -- 2885834784
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ff17dc24" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"536d2720"; -- 1399662368
        operand2 <= x"acee83a2"; -- 2901312418
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffefa7a2" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"df63ab6f"; -- 3747851119
        operand2 <= x"2b78e210"; -- 729342480
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ff7beb7f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f01dc0af"; -- 4028481711
        operand2 <= x"229cebfa"; -- 580709370
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f29debff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3d586fd0"; -- 1029205968
        operand2 <= x"3d0e1532"; -- 1024333106
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3d5e7ff2" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e9f4f360"; -- 3925144416
        operand2 <= x"5b46c5d6"; -- 1531364822
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fbf6f7f6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9b56567f"; -- 2606126719
        operand2 <= x"081072d9"; -- 135295705
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9b5676ff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d7a91936"; -- 3618183478
        operand2 <= x"020aa055"; -- 34250837
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d7abb977" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dc06420f"; -- 3691397647
        operand2 <= x"1fc1b6b5"; -- 532788917
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"dfc7f6bf" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b6c50c4f"; -- 3066367055
        operand2 <= x"622886e2"; -- 1646823138
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f6ed8eef" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"da9728df"; -- 3667339487
        operand2 <= x"17b78f01"; -- 397905665
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"dfb7afdf" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bb8fcaa4"; -- 3146762916
        operand2 <= x"860c8072"; -- 2248966258
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bf8fcaf6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"cefddca9"; -- 3472743593
        operand2 <= x"0c74f391"; -- 208991121
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"cefdffb9" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0f2d8321"; -- 254640929
        operand2 <= x"61f510d8"; -- 1643450584
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6ffd93f9" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3be01a2b"; -- 1004542507
        operand2 <= x"227f6b9b"; -- 578775963
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3bff7bbb" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6afb6161"; -- 1794859361
        operand2 <= x"ec1a0571"; -- 3961128305
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"eefb6571" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"79275f66"; -- 2032623462
        operand2 <= x"28106841"; -- 672163905
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"79377f67" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b7657f71"; -- 3076882289
        operand2 <= x"e8da40ef"; -- 3906617583
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffff7fff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ef09ecef"; -- 4010405103
        operand2 <= x"cde59b09"; -- 3454376713
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"efedffef" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c3c976f8"; -- 3284760312
        operand2 <= x"46418c28"; -- 1178700840
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c7c9fef8" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"437fc214"; -- 1132446228
        operand2 <= x"33f597b5"; -- 871733173
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"73ffd7b5" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"eb30c21c"; -- 3945841180
        operand2 <= x"605181a1"; -- 1615954337
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"eb71c3bd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2762214c"; -- 660742476
        operand2 <= x"1f4f80d5"; -- 525304021
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3f6fa1dd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2a30874e"; -- 707823438
        operand2 <= x"608c8d1c"; -- 1619823900
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6abc8f5e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fae469ce"; -- 4209273294
        operand2 <= x"80db6f18"; -- 2161864472
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"faff6fde" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0e9384d9"; -- 244548825
        operand2 <= x"8105613a"; -- 2164613434
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8f97e5fb" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1f739c1d"; -- 527670301
        operand2 <= x"c873606a"; -- 3363004522
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"df73fc7f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"79b5c492"; -- 2041955474
        operand2 <= x"d34a8134"; -- 3544875316
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fbffc5b6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2520477e"; -- 622872446
        operand2 <= x"bb537ae5"; -- 3142810341
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bf737fff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6291c066"; -- 1653719142
        operand2 <= x"f8abb130"; -- 4172001584
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fabbf176" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b81fd653"; -- 3089094227
        operand2 <= x"0a74f982"; -- 175438210
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ba7fffd3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"cd9e39b9"; -- 3449698745
        operand2 <= x"db60d095"; -- 3680555157
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"dffef9bd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4a94f8d2"; -- 1251277010
        operand2 <= x"3187b761"; -- 830977889
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7b97fff3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"acf8715f"; -- 2901963103
        operand2 <= x"eaac6b42"; -- 3937168194
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"eefc7b5f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"47a50977"; -- 1201998199
        operand2 <= x"c6f33c81"; -- 3337829505
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c7f73df7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f45160b4"; -- 4098973876
        operand2 <= x"3e8de5cc"; -- 1049486796
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fedde5fc" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7ff7061a"; -- 2146895386
        operand2 <= x"62c8ef0f"; -- 1657335567
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7fffef1f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dff249f1"; -- 3757197809
        operand2 <= x"a89cb945"; -- 2828843333
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fffef9f5" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"820c0db1"; -- 2181828017
        operand2 <= x"70af256a"; -- 1890526570
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f2af2dfb" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8d3d0226"; -- 2369585702
        operand2 <= x"1e53f871"; -- 508819569
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9f7ffa77" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"727a8563"; -- 1920632163
        operand2 <= x"86d62c3e"; -- 2262182974
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f6fead7f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ce56ac8d"; -- 3461786765
        operand2 <= x"6bc1f634"; -- 1807873588
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"efd7febd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"11cc77e9"; -- 298612713
        operand2 <= x"6b021540"; -- 1795298624
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7bce77e9" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"418c8033"; -- 1099726899
        operand2 <= x"5f45e4a1"; -- 1598416033
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"5fcde4b3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ab72bb8c"; -- 2876423052
        operand2 <= x"0b0c19cc"; -- 185342412
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ab7ebbcc" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1fc1b3b1"; -- 532788145
        operand2 <= x"8829eabf"; -- 2284448447
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9fe9fbbf" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2a7fecec"; -- 713026796
        operand2 <= x"63bc87f9"; -- 1673299961
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6bffeffd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2644dc06"; -- 642046982
        operand2 <= x"360d8661"; -- 906856033
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"364dde67" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dfcdbe31"; -- 3754802737
        operand2 <= x"4a279dae"; -- 1244110254
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"dfefbfbf" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b7402dcc"; -- 3074436556
        operand2 <= x"0fed2fd3"; -- 267202515
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bfed2fdf" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"42574085"; -- 1113014405
        operand2 <= x"a8771481"; -- 2826376321
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ea775485" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bd9766b4"; -- 3180816052
        operand2 <= x"78fab464"; -- 2029696100
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fdfff6f4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"cfa7a72a"; -- 3483871018
        operand2 <= x"5a335977"; -- 1513314679
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"dfb7ff7f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"854abb8f"; -- 2236267407
        operand2 <= x"8c53fe9d"; -- 2354314909
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8d5bff9f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a779d638"; -- 2809779768
        operand2 <= x"e56f8934"; -- 3849292084
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"e77fdf3c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1dfbc4a5"; -- 503039141
        operand2 <= x"60b11aea"; -- 1622219498
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7dfbdeef" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2f162508"; -- 789980424
        operand2 <= x"9f3654fa"; -- 2671138042
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bf3675fa" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c719a8c3"; -- 3340347587
        operand2 <= x"fe61ceb6"; -- 4267822774
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ff79eef7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a85559e9"; -- 2824165865
        operand2 <= x"ad81a29e"; -- 2910954142
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"add5fbff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3b918f72"; -- 999395186
        operand2 <= x"ec3efe5d"; -- 3963551325
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffbfff7f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0f4e3bee"; -- 256785390
        operand2 <= x"64258d8f"; -- 1680182671
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6f6fbfef" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fcf14ccd"; -- 4243672269
        operand2 <= x"41c38981"; -- 1103333761
        ALUOp <= "001";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fdf3cdcd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2137bb8c"; -- 557300620
        operand2 <= x"f04fbbb3"; -- 4031757235
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d178003f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"73e1d94a"; -- 1944181066
        operand2 <= x"eac6c772"; -- 3938895730
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"99271e38" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ec8e6bc8"; -- 3968756680
        operand2 <= x"af42bfae"; -- 2940387246
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"43ccd466" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2fc468ef"; -- 801401071
        operand2 <= x"df7b27a4"; -- 3749390244
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f0bf4f4b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8c73cbe8"; -- 2356399080
        operand2 <= x"33af33cc"; -- 867120076
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bfdcf824" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1fdd9797"; -- 534615959
        operand2 <= x"a450e9d3"; -- 2756766163
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bb8d7e44" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7cfe77f3"; -- 2097051635
        operand2 <= x"b21514b2"; -- 2987726002
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ceeb6341" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"38e0d5cd"; -- 954258893
        operand2 <= x"edfce08a"; -- 3992772746
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d51c3547" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b1f6568e"; -- 2985711246
        operand2 <= x"1c7b9f9c"; -- 477863836
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ad8dc912" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c48dde4a"; -- 3297631818
        operand2 <= x"075db4c6"; -- 123581638
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c3d06a8c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"20a0c788"; -- 547407752
        operand2 <= x"6792e99f"; -- 1737681311
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"47322e17" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f60dedde"; -- 4128107998
        operand2 <= x"a7609d2b"; -- 2808126763
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"516d70f5" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"67220b4f"; -- 1730284367
        operand2 <= x"5f40de45"; -- 1598086725
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3862d50a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"529525ad"; -- 1385506221
        operand2 <= x"932afcc3"; -- 2469067971
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c1bfd96e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4e9709b2"; -- 1318521266
        operand2 <= x"67264048"; -- 1730560072
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"29b149fa" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dec2a838"; -- 3737299000
        operand2 <= x"1d1fe185"; -- 488628613
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c3dd49bd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"97aa1405"; -- 2544505861
        operand2 <= x"d1efa5d2"; -- 3522143698
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4645b1d7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4094efa2"; -- 1083502498
        operand2 <= x"86b49c8f"; -- 2259983503
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c620732d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"92fb691d"; -- 2465949981
        operand2 <= x"8ed74ff7"; -- 2396475383
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1c2c26ea" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ff3b66f3"; -- 4282083059
        operand2 <= x"ea072eae"; -- 3926339246
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"153c485d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"810333da"; -- 2164470746
        operand2 <= x"63009083"; -- 1660981379
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"e203a359" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6cf419be"; -- 1827936702
        operand2 <= x"ef47c556"; -- 4014458198
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"83b3dce8" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d889e2c5"; -- 3632915141
        operand2 <= x"c0b82626"; -- 3233293862
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1831c4e3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"936786c8"; -- 2473035464
        operand2 <= x"7d2c0ad7"; -- 2100038359
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ee4b8c1f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"19e56e4f"; -- 434466383
        operand2 <= x"aa46c385"; -- 2856764293
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b3a3adca" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"41ca71a0"; -- 1103786400
        operand2 <= x"d0b53a10"; -- 3501537808
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"917f4bb0" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1be336c1"; -- 467875521
        operand2 <= x"a43fc934"; -- 2755643700
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bfdcfff5" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"84a2aeef"; -- 2225254127
        operand2 <= x"81dce945"; -- 2178738501
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"057e47aa" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b9d76ced"; -- 3117903085
        operand2 <= x"2f0d6dcb"; -- 789409227
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"96da0126" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"53316d99"; -- 1395748249
        operand2 <= x"e3cc4c43"; -- 3821816899
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b0fd21da" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6097a6b4"; -- 1620551348
        operand2 <= x"f8a23832"; -- 4171380786
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"98359e86" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e2f7e4fe"; -- 3807896830
        operand2 <= x"c7c709b2"; -- 3351710130
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2530ed4c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a422dbcf"; -- 2753747919
        operand2 <= x"973f85e3"; -- 2537522659
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"331d5e2c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"57068e30"; -- 1460047408
        operand2 <= x"ddc413b7"; -- 3720614839
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8ac29d87" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3d3c25d2"; -- 1027352018
        operand2 <= x"3b5a18be"; -- 995760318
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"06663d6c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c2973c77"; -- 3264691319
        operand2 <= x"0a7c1e7b"; -- 175906427
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c8eb220c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a30725ae"; -- 2735154606
        operand2 <= x"a8a5e670"; -- 2829444720
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0ba2c3de" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"cb575ae2"; -- 3411499746
        operand2 <= x"33bd6277"; -- 868049527
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f8ea3895" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"119cfeca"; -- 295501514
        operand2 <= x"5b051d42"; -- 1527061826
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4a99e388" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4a3935bc"; -- 1245263292
        operand2 <= x"9eb18fbf"; -- 2662436799
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d488ba03" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bd8426e1"; -- 3179554529
        operand2 <= x"546c5b81"; -- 1416387457
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"e9e87d60" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"cd015b3d"; -- 3439418173
        operand2 <= x"91abcf8b"; -- 2443956107
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"5caa94b6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5eaa2869"; -- 1588209769
        operand2 <= x"4304dae6"; -- 1124391654
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1daef28f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"06c617db"; -- 113645531
        operand2 <= x"bf64fa25"; -- 3211065893
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b9a2edfe" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c0ff85c4"; -- 3237971396
        operand2 <= x"7de042a8"; -- 2111849128
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bd1fc76c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d45251b8"; -- 3562164664
        operand2 <= x"a446d07f"; -- 2756104319
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"701481c7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"88b55173"; -- 2293584243
        operand2 <= x"39c6ca05"; -- 969329157
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b1739b76" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7de91510"; -- 2112427280
        operand2 <= x"95f4c5bd"; -- 2515846589
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"e81dd0ad" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"45400d38"; -- 1161825592
        operand2 <= x"e2e1a8a1"; -- 3806439585
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a7a1a599" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"798d2729"; -- 2039293737
        operand2 <= x"f2252628"; -- 4062520872
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8ba80101" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"94498418"; -- 2487845912
        operand2 <= x"b29ecf8d"; -- 2996752269
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"26d74b95" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3c9321b6"; -- 1016275382
        operand2 <= x"6e5756ff"; -- 1851217663
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"52c47749" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"11374c88"; -- 288836744
        operand2 <= x"7293683c"; -- 1922263100
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"63a424b4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8a519db3"; -- 2320604595
        operand2 <= x"724cb1e3"; -- 1917628899
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f81d2c50" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"85d466e4"; -- 2245289700
        operand2 <= x"9cf0fd09"; -- 2633039113
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"19249bed" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d8c8a4c0"; -- 3637028032
        operand2 <= x"91d3bca6"; -- 2446572710
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"491b1866" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a04f0ee1"; -- 2689535713
        operand2 <= x"850e6940"; -- 2232314176
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"254167a1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b1fe2fac"; -- 2986225580
        operand2 <= x"ef9f5500"; -- 4020196608
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"5e617aac" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6545a642"; -- 1699063362
        operand2 <= x"c053c5c6"; -- 3226715590
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a5166384" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"da260fd5"; -- 3659927509
        operand2 <= x"beef8de7"; -- 3203370471
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"64c98232" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"710b2b40"; -- 1896557376
        operand2 <= x"6bc14ed1"; -- 1807830737
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1aca6591" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"50874ae1"; -- 1351043809
        operand2 <= x"7dec83bd"; -- 2112652221
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2d6bc95c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2edfc955"; -- 786418005
        operand2 <= x"115074c7"; -- 290485447
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3f8fbd92" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6bc88202"; -- 1808302594
        operand2 <= x"d80dc32e"; -- 3624780590
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b3c5412c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"844d6f5e"; -- 2219667294
        operand2 <= x"60074262"; -- 1611088482
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"e44a2d3c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"246008dd"; -- 610273501
        operand2 <= x"156a798c"; -- 359299468
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"310a7151" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1f3080fb"; -- 523272443
        operand2 <= x"ca54fe01"; -- 3394567681
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d5647efa" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0d08a393"; -- 218669971
        operand2 <= x"6e3d2025"; -- 1849499685
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"633583b6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4bd281c8"; -- 1272086984
        operand2 <= x"1d27e47c"; -- 489153660
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"56f565b4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9e1e90e4"; -- 2652803300
        operand2 <= x"ec105642"; -- 3960493634
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"720ec6a6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5c9f927a"; -- 1553961594
        operand2 <= x"8dde1c61"; -- 2380143713
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d1418e1b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6bc5e8ac"; -- 1808132268
        operand2 <= x"01e24a3a"; -- 31607354
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6a27a296" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dd78940a"; -- 3715666954
        operand2 <= x"77cdd78c"; -- 2009978764
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"aab54386" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f49b3dfa"; -- 4103814650
        operand2 <= x"ffb0a2e6"; -- 4289766118
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0b2b9f1c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"427a75af"; -- 1115321775
        operand2 <= x"ecefa834"; -- 3975129140
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ae95dd9b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f8a40d1e"; -- 4171500830
        operand2 <= x"5fbe903a"; -- 1606324282
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a71a9d24" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a3d798d7"; -- 2748815575
        operand2 <= x"bd810ed4"; -- 3179351764
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1e569603" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"06b0c382"; -- 112247682
        operand2 <= x"961180ed"; -- 2517729517
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"90a1436f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a751be65"; -- 2807152229
        operand2 <= x"39084bb7"; -- 956844983
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9e59f5d2" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"821e2f6d"; -- 2183016301
        operand2 <= x"05738bde"; -- 91458526
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"876da4b3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e5c2e551"; -- 3854755153
        operand2 <= x"5027795f"; -- 1344764255
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b5e59c0e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"23baa488"; -- 599434376
        operand2 <= x"db3eeead"; -- 3678334637
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f8844a25" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0f5c0768"; -- 257689448
        operand2 <= x"85f10d24"; -- 2247167268
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8aad0a4c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5820e265"; -- 1478550117
        operand2 <= x"6008bcf3"; -- 1611185395
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"38285e96" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2d8e013e"; -- 764281150
        operand2 <= x"05b27f38"; -- 95584056
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"283c7e06" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2111c78e"; -- 554813326
        operand2 <= x"dd524227"; -- 3713155623
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fc4385a9" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c15d923c"; -- 3244134972
        operand2 <= x"56a50d06"; -- 1453657350
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"97f89f3a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"115beb85"; -- 291236741
        operand2 <= x"79e4b095"; -- 2045030549
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"68bf5b10" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3c1f2120"; -- 1008673056
        operand2 <= x"1a6b84da"; -- 443253978
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2674a5fa" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9ee5d8b3"; -- 2665863347
        operand2 <= x"977f10f3"; -- 2541687027
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"099ac840" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"aee4e665"; -- 2934236773
        operand2 <= x"51a0437f"; -- 1369457535
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ff44a51a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dc982806"; -- 3700959238
        operand2 <= x"127d9451"; -- 310219857
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"cee5bc57" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"de1c7c72"; -- 3726408818
        operand2 <= x"8bf3eaa9"; -- 2348018345
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"55ef96db" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5decebe4"; -- 1575807972
        operand2 <= x"e35e2f25"; -- 3814600485
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"beb2c4c1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c4fc96b1"; -- 3304887985
        operand2 <= x"23e228a7"; -- 602024103
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"e71ebe16" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0b000121"; -- 184549665
        operand2 <= x"33784634"; -- 863520308
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"38784715" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"04198927"; -- 68782375
        operand2 <= x"f5ff20b9"; -- 4127137977
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f1e6a99e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"32d96b1b"; -- 853109531
        operand2 <= x"9cef659b"; -- 2632934811
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ae360e80" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b473a6c6"; -- 3027478214
        operand2 <= x"fa645c96"; -- 4200881302
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4e17fa50" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"88b360bd"; -- 2293457085
        operand2 <= x"f5169808"; -- 4111898632
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7da5f8b5" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"59b335ee"; -- 1504916974
        operand2 <= x"a219a2ba"; -- 2719589050
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fbaa9754" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"cd3f4a92"; -- 3443477138
        operand2 <= x"c985ea35"; -- 3380996661
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"04baa0a7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bbefb67b"; -- 3153049211
        operand2 <= x"ae3807b7"; -- 2922907575
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"15d7b1cc" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bbd3b499"; -- 3151213721
        operand2 <= x"21d2a01b"; -- 567451675
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9a011482" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c5b8e5a1"; -- 3317228961
        operand2 <= x"ff3f43bd"; -- 4282336189
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3a87a61c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"22bce20c"; -- 582803980
        operand2 <= x"26ba4271"; -- 649740913
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0406a07d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ed0fc07f"; -- 3977232511
        operand2 <= x"d4089da0"; -- 3557334432
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"39075ddf" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dd8edd20"; -- 3717127456
        operand2 <= x"5ba25370"; -- 1537364848
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"862c8e50" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"58480255"; -- 1481114197
        operand2 <= x"2510f73f"; -- 621868863
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7d58f56a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ee22b293"; -- 3995251347
        operand2 <= x"f70879f6"; -- 4144527862
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"192acb65" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"45f86c3f"; -- 1173908543
        operand2 <= x"cbf20c99"; -- 3421637785
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8e0a60a6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0368573b"; -- 57169723
        operand2 <= x"79ebc56e"; -- 2045494638
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7a839255" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7b27588d"; -- 2066176141
        operand2 <= x"15e8b820"; -- 367573024
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6ecfe0ad" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"97e67208"; -- 2548462088
        operand2 <= x"729a55b5"; -- 1922717109
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"e57c27bd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"34f1cda4"; -- 888262052
        operand2 <= x"a29629b0"; -- 2727750064
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9667e414" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"01f2e928"; -- 32696616
        operand2 <= x"6385e3a2"; -- 1669718946
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"62770a8a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"88745e2d"; -- 2289327661
        operand2 <= x"ea584a76"; -- 3931654774
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"622c145b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a6764142"; -- 2792767810
        operand2 <= x"7ed6ec69"; -- 2128014441
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d8a0ad2b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8158a33f"; -- 2170069823
        operand2 <= x"e5915c8e"; -- 3851508878
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"64c9ffb1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"830df103"; -- 2198728963
        operand2 <= x"cefafa65"; -- 3472554597
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4df70b66" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4b94b875"; -- 1268037749
        operand2 <= x"e458cb7f"; -- 3831024511
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"afcc730a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4e308e0a"; -- 1311804938
        operand2 <= x"74610c57"; -- 1952517207
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3a51825d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"36bca71a"; -- 918333210
        operand2 <= x"15353b23"; -- 355810083
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"23899c39" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fed9b287"; -- 4275679879
        operand2 <= x"fc56c860"; -- 4233545824
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"028f7ae7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"07efb355"; -- 133149525
        operand2 <= x"9543759f"; -- 2504226207
        ALUOp <= "010";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"92acc6ca" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9e905b21"; -- 2660260641
        operand2 <= x"8acabfd0"; -- 2328543184
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9e905b21"; -- 2660260641
        operand2 <= x"8acabfd0"; -- 2328543184
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"aace1662"; -- 2865632866
        operand2 <= x"186bdc27"; -- 409721895
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"aace1662"; -- 2865632866
        operand2 <= x"186bdc27"; -- 409721895
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ee6bee0c"; -- 4000050700
        operand2 <= x"b98ba121"; -- 3112935713
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ee6bee0c"; -- 4000050700
        operand2 <= x"b98ba121"; -- 3112935713
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d05f0eef"; -- 3495890671
        operand2 <= x"b18f20af"; -- 2978947247
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d05f0eef"; -- 3495890671
        operand2 <= x"b18f20af"; -- 2978947247
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3c071477"; -- 1007096951
        operand2 <= x"2ad21166"; -- 718410086
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3c071477"; -- 1007096951
        operand2 <= x"2ad21166"; -- 718410086
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9751541e"; -- 2538689566
        operand2 <= x"674de064"; -- 1733156964
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9751541e"; -- 2538689566
        operand2 <= x"674de064"; -- 1733156964
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2c0e9156"; -- 739152214
        operand2 <= x"5b33715e"; -- 1530098014
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2c0e9156"; -- 739152214
        operand2 <= x"5b33715e"; -- 1530098014
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8f770d73"; -- 2406944115
        operand2 <= x"79b7a47b"; -- 2042078331
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8f770d73"; -- 2406944115
        operand2 <= x"79b7a47b"; -- 2042078331
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ae8dddfd"; -- 2928532989
        operand2 <= x"b150afb2"; -- 2974855090
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ae8dddfd"; -- 2928532989
        operand2 <= x"b150afb2"; -- 2974855090
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"adf1f381"; -- 2918314881
        operand2 <= x"12bdd57f"; -- 314430847
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"adf1f381"; -- 2918314881
        operand2 <= x"12bdd57f"; -- 314430847
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"65a035fc"; -- 1704998396
        operand2 <= x"5c6ecad9"; -- 1550764761
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"65a035fc"; -- 1704998396
        operand2 <= x"5c6ecad9"; -- 1550764761
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7af54665"; -- 2062894693
        operand2 <= x"1e32cac3"; -- 506645187
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7af54665"; -- 2062894693
        operand2 <= x"1e32cac3"; -- 506645187
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9a255d48"; -- 2586139976
        operand2 <= x"e5ecc300"; -- 3857498880
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9a255d48"; -- 2586139976
        operand2 <= x"e5ecc300"; -- 3857498880
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"14de2698"; -- 350103192
        operand2 <= x"f9f75204"; -- 4193735172
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"14de2698"; -- 350103192
        operand2 <= x"f9f75204"; -- 4193735172
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c121c2df"; -- 3240215263
        operand2 <= x"4cc4ecd3"; -- 1287974099
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c121c2df"; -- 3240215263
        operand2 <= x"4cc4ecd3"; -- 1287974099
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"919279da"; -- 2442295770
        operand2 <= x"301bc85b"; -- 807127131
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"919279da"; -- 2442295770
        operand2 <= x"301bc85b"; -- 807127131
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"96463dca"; -- 2521185738
        operand2 <= x"e201e6f3"; -- 3791775475
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"96463dca"; -- 2521185738
        operand2 <= x"e201e6f3"; -- 3791775475
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"331bb9d5"; -- 857455061
        operand2 <= x"1c425a58"; -- 474110552
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"331bb9d5"; -- 857455061
        operand2 <= x"1c425a58"; -- 474110552
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"69545471"; -- 1767134321
        operand2 <= x"55bb2b88"; -- 1438329736
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"69545471"; -- 1767134321
        operand2 <= x"55bb2b88"; -- 1438329736
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"90447d4c"; -- 2420407628
        operand2 <= x"e4140496"; -- 3826517142
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"90447d4c"; -- 2420407628
        operand2 <= x"e4140496"; -- 3826517142
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7363df9c"; -- 1935925148
        operand2 <= x"0f6dfd3b"; -- 258866491
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7363df9c"; -- 1935925148
        operand2 <= x"0f6dfd3b"; -- 258866491
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1f640033"; -- 526647347
        operand2 <= x"2d5b9362"; -- 760976226
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1f640033"; -- 526647347
        operand2 <= x"2d5b9362"; -- 760976226
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"431ca5ed"; -- 1125950957
        operand2 <= x"befd8453"; -- 3204285523
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"431ca5ed"; -- 1125950957
        operand2 <= x"befd8453"; -- 3204285523
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"35dd661c"; -- 903702044
        operand2 <= x"b601035e"; -- 3053519710
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"35dd661c"; -- 903702044
        operand2 <= x"b601035e"; -- 3053519710
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"55505801"; -- 1431328769
        operand2 <= x"16f5202d"; -- 385163309
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"55505801"; -- 1431328769
        operand2 <= x"16f5202d"; -- 385163309
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1a0aa863"; -- 436906083
        operand2 <= x"d6ee3fa2"; -- 3605938082
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1a0aa863"; -- 436906083
        operand2 <= x"d6ee3fa2"; -- 3605938082
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8f8cd7f4"; -- 2408372212
        operand2 <= x"d5d5b661"; -- 3587552865
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8f8cd7f4"; -- 2408372212
        operand2 <= x"d5d5b661"; -- 3587552865
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"14e1a121"; -- 350331169
        operand2 <= x"1efdf818"; -- 519960600
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"14e1a121"; -- 350331169
        operand2 <= x"1efdf818"; -- 519960600
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ed6f28f3"; -- 3983485171
        operand2 <= x"61555246"; -- 1632981574
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ed6f28f3"; -- 3983485171
        operand2 <= x"61555246"; -- 1632981574
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6d030e93"; -- 1828916883
        operand2 <= x"7f863545"; -- 2139501893
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6d030e93"; -- 1828916883
        operand2 <= x"7f863545"; -- 2139501893
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"803bc2db"; -- 2151400155
        operand2 <= x"89827ab2"; -- 2307029682
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"803bc2db"; -- 2151400155
        operand2 <= x"89827ab2"; -- 2307029682
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e20d009e"; -- 3792502942
        operand2 <= x"9d796361"; -- 2641978209
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e20d009e"; -- 3792502942
        operand2 <= x"9d796361"; -- 2641978209
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0c2e7378"; -- 204370808
        operand2 <= x"69617a46"; -- 1767995974
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0c2e7378"; -- 204370808
        operand2 <= x"69617a46"; -- 1767995974
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9ca0c183"; -- 2627780995
        operand2 <= x"bab1ea9f"; -- 3132222111
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9ca0c183"; -- 2627780995
        operand2 <= x"bab1ea9f"; -- 3132222111
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7e818869"; -- 2122418281
        operand2 <= x"345a41e2"; -- 878330338
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7e818869"; -- 2122418281
        operand2 <= x"345a41e2"; -- 878330338
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1f07e9ec"; -- 520612332
        operand2 <= x"8ebeda07"; -- 2394872327
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1f07e9ec"; -- 520612332
        operand2 <= x"8ebeda07"; -- 2394872327
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5964c9f7"; -- 1499777527
        operand2 <= x"eb3b9a85"; -- 3946551941
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5964c9f7"; -- 1499777527
        operand2 <= x"eb3b9a85"; -- 3946551941
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"02bd199c"; -- 45947292
        operand2 <= x"e5418e8f"; -- 3846278799
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"02bd199c"; -- 45947292
        operand2 <= x"e5418e8f"; -- 3846278799
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e464783b"; -- 3831789627
        operand2 <= x"f63fff05"; -- 4131389189
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e464783b"; -- 3831789627
        operand2 <= x"f63fff05"; -- 4131389189
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"aeffb228"; -- 2935992872
        operand2 <= x"7985326d"; -- 2038772333
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"aeffb228"; -- 2935992872
        operand2 <= x"7985326d"; -- 2038772333
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"211ba55c"; -- 555459932
        operand2 <= x"a65f2e2a"; -- 2791255594
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"211ba55c"; -- 555459932
        operand2 <= x"a65f2e2a"; -- 2791255594
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"227564a6"; -- 578118822
        operand2 <= x"c6c62575"; -- 3334874485
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"227564a6"; -- 578118822
        operand2 <= x"c6c62575"; -- 3334874485
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4fca39cf"; -- 1338653135
        operand2 <= x"de7d4d03"; -- 3732753667
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4fca39cf"; -- 1338653135
        operand2 <= x"de7d4d03"; -- 3732753667
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ab3f5351"; -- 2873054033
        operand2 <= x"9652ea2e"; -- 2522016302
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ab3f5351"; -- 2873054033
        operand2 <= x"9652ea2e"; -- 2522016302
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"29f691c4"; -- 704025028
        operand2 <= x"d26dadc0"; -- 3530403264
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"29f691c4"; -- 704025028
        operand2 <= x"d26dadc0"; -- 3530403264
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5a15661e"; -- 1511351838
        operand2 <= x"7e32e992"; -- 2117265810
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5a15661e"; -- 1511351838
        operand2 <= x"7e32e992"; -- 2117265810
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"40ea6eba"; -- 1089105594
        operand2 <= x"5c3c9aef"; -- 1547475695
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"40ea6eba"; -- 1089105594
        operand2 <= x"5c3c9aef"; -- 1547475695
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"70f15b44"; -- 1894865732
        operand2 <= x"0cd8399f"; -- 215497119
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"70f15b44"; -- 1894865732
        operand2 <= x"0cd8399f"; -- 215497119
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"45b40165"; -- 1169424741
        operand2 <= x"a5c52b04"; -- 2781162244
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"45b40165"; -- 1169424741
        operand2 <= x"a5c52b04"; -- 2781162244
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b66bcaee"; -- 3060517614
        operand2 <= x"4c94e1bd"; -- 1284825533
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b66bcaee"; -- 3060517614
        operand2 <= x"4c94e1bd"; -- 1284825533
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3618d3d6"; -- 907596758
        operand2 <= x"6360670c"; -- 1667262220
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3618d3d6"; -- 907596758
        operand2 <= x"6360670c"; -- 1667262220
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d5409e06"; -- 3577781766
        operand2 <= x"9ca8b025"; -- 2628300837
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d5409e06"; -- 3577781766
        operand2 <= x"9ca8b025"; -- 2628300837
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6045fd92"; -- 1615199634
        operand2 <= x"1bfca97e"; -- 469543294
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6045fd92"; -- 1615199634
        operand2 <= x"1bfca97e"; -- 469543294
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1483eedd"; -- 344190685
        operand2 <= x"3f603a37"; -- 1063270967
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1483eedd"; -- 344190685
        operand2 <= x"3f603a37"; -- 1063270967
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9435e3fd"; -- 2486559741
        operand2 <= x"6a5b726d"; -- 1784377965
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9435e3fd"; -- 2486559741
        operand2 <= x"6a5b726d"; -- 1784377965
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b329a474"; -- 3005850740
        operand2 <= x"b56e5308"; -- 3043906312
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b329a474"; -- 3005850740
        operand2 <= x"b56e5308"; -- 3043906312
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e3c631e6"; -- 3821416934
        operand2 <= x"98ba2e26"; -- 2562338342
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e3c631e6"; -- 3821416934
        operand2 <= x"98ba2e26"; -- 2562338342
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e6363f1d"; -- 3862314781
        operand2 <= x"3834421e"; -- 942948894
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e6363f1d"; -- 3862314781
        operand2 <= x"3834421e"; -- 942948894
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2c239ca8"; -- 740531368
        operand2 <= x"0902ad43"; -- 151170371
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2c239ca8"; -- 740531368
        operand2 <= x"0902ad43"; -- 151170371
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"99d08872"; -- 2580580466
        operand2 <= x"070baae1"; -- 118205153
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"99d08872"; -- 2580580466
        operand2 <= x"070baae1"; -- 118205153
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0529f705"; -- 86636293
        operand2 <= x"02d944d0"; -- 47793360
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0529f705"; -- 86636293
        operand2 <= x"02d944d0"; -- 47793360
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fc6ef0b0"; -- 4235129008
        operand2 <= x"ccf17452"; -- 3438376018
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fc6ef0b0"; -- 4235129008
        operand2 <= x"ccf17452"; -- 3438376018
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2203ce28"; -- 570674728
        operand2 <= x"2ffd6019"; -- 805134361
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2203ce28"; -- 570674728
        operand2 <= x"2ffd6019"; -- 805134361
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a284c19b"; -- 2726609307
        operand2 <= x"0f5402ae"; -- 257163950
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a284c19b"; -- 2726609307
        operand2 <= x"0f5402ae"; -- 257163950
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7e9524ea"; -- 2123703530
        operand2 <= x"84b01787"; -- 2226132871
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7e9524ea"; -- 2123703530
        operand2 <= x"84b01787"; -- 2226132871
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6502ff57"; -- 1694695255
        operand2 <= x"d5169b8d"; -- 3575028621
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6502ff57"; -- 1694695255
        operand2 <= x"d5169b8d"; -- 3575028621
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f475d928"; -- 4101364008
        operand2 <= x"0f313620"; -- 254883360
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f475d928"; -- 4101364008
        operand2 <= x"0f313620"; -- 254883360
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a83758ef"; -- 2822199535
        operand2 <= x"7b19de6e"; -- 2065292910
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a83758ef"; -- 2822199535
        operand2 <= x"7b19de6e"; -- 2065292910
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"88dac702"; -- 2296039170
        operand2 <= x"470c43e2"; -- 1191986146
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"88dac702"; -- 2296039170
        operand2 <= x"470c43e2"; -- 1191986146
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e8ca433c"; -- 3905569596
        operand2 <= x"7a1d0617"; -- 2048722455
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e8ca433c"; -- 3905569596
        operand2 <= x"7a1d0617"; -- 2048722455
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9b02e2db"; -- 2600657627
        operand2 <= x"81bffc03"; -- 2176842755
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9b02e2db"; -- 2600657627
        operand2 <= x"81bffc03"; -- 2176842755
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"abafecf5"; -- 2880433397
        operand2 <= x"733e27c4"; -- 1933453252
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"abafecf5"; -- 2880433397
        operand2 <= x"733e27c4"; -- 1933453252
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c7936fcd"; -- 3348328397
        operand2 <= x"bb0bad57"; -- 3138104663
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c7936fcd"; -- 3348328397
        operand2 <= x"bb0bad57"; -- 3138104663
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c98eecad"; -- 3381587117
        operand2 <= x"0d3dd6b2"; -- 222156466
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c98eecad"; -- 3381587117
        operand2 <= x"0d3dd6b2"; -- 222156466
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"53fb2664"; -- 1408968292
        operand2 <= x"b5e773b9"; -- 3051844537
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"53fb2664"; -- 1408968292
        operand2 <= x"b5e773b9"; -- 3051844537
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b1e615bb"; -- 2984646075
        operand2 <= x"3b3a87ec"; -- 993691628
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b1e615bb"; -- 2984646075
        operand2 <= x"3b3a87ec"; -- 993691628
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9612b4a2"; -- 2517808290
        operand2 <= x"d329871a"; -- 3542714138
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9612b4a2"; -- 2517808290
        operand2 <= x"d329871a"; -- 3542714138
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"251dd478"; -- 622711928
        operand2 <= x"e4129583"; -- 3826423171
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"251dd478"; -- 622711928
        operand2 <= x"e4129583"; -- 3826423171
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1c7b9002"; -- 477859842
        operand2 <= x"47e95563"; -- 1206474083
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1c7b9002"; -- 477859842
        operand2 <= x"47e95563"; -- 1206474083
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0f3df496"; -- 255718550
        operand2 <= x"36c973b1"; -- 919172017
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0f3df496"; -- 255718550
        operand2 <= x"36c973b1"; -- 919172017
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"cf30dbc4"; -- 3476085700
        operand2 <= x"8decaef9"; -- 2381098745
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"cf30dbc4"; -- 3476085700
        operand2 <= x"8decaef9"; -- 2381098745
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fcc85931"; -- 4240988465
        operand2 <= x"3bd553bd"; -- 1003836349
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fcc85931"; -- 4240988465
        operand2 <= x"3bd553bd"; -- 1003836349
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"46d1f4e1"; -- 1188164833
        operand2 <= x"af4b25ef"; -- 2940937711
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"46d1f4e1"; -- 1188164833
        operand2 <= x"af4b25ef"; -- 2940937711
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bfaa68d0"; -- 3215616208
        operand2 <= x"8d14b97b"; -- 2366945659
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bfaa68d0"; -- 3215616208
        operand2 <= x"8d14b97b"; -- 2366945659
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"413b7f5d"; -- 1094418269
        operand2 <= x"8b928aec"; -- 2341636844
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"413b7f5d"; -- 1094418269
        operand2 <= x"8b928aec"; -- 2341636844
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"031fcbb2"; -- 52415410
        operand2 <= x"6347400a"; -- 1665613834
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"031fcbb2"; -- 52415410
        operand2 <= x"6347400a"; -- 1665613834
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0c93c1b5"; -- 211009973
        operand2 <= x"41eb9557"; -- 1105958231
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0c93c1b5"; -- 211009973
        operand2 <= x"41eb9557"; -- 1105958231
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3aeaefde"; -- 988475358
        operand2 <= x"061dc960"; -- 102615392
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3aeaefde"; -- 988475358
        operand2 <= x"061dc960"; -- 102615392
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d5fbbbad"; -- 3590044589
        operand2 <= x"f1a10d8b"; -- 4053863819
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d5fbbbad"; -- 3590044589
        operand2 <= x"f1a10d8b"; -- 4053863819
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3684dc4a"; -- 914676810
        operand2 <= x"f5fdf950"; -- 4127062352
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3684dc4a"; -- 914676810
        operand2 <= x"f5fdf950"; -- 4127062352
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ba8e84ee"; -- 3129902318
        operand2 <= x"9c72cadc"; -- 2624768732
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ba8e84ee"; -- 3129902318
        operand2 <= x"9c72cadc"; -- 2624768732
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"158737dc"; -- 361183196
        operand2 <= x"5b047a3a"; -- 1527020090
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"158737dc"; -- 361183196
        operand2 <= x"5b047a3a"; -- 1527020090
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e5e7dcbb"; -- 3857177787
        operand2 <= x"a67110c7"; -- 2792427719
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e5e7dcbb"; -- 3857177787
        operand2 <= x"a67110c7"; -- 2792427719
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a2eff83b"; -- 2733635643
        operand2 <= x"348cadd9"; -- 881634777
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a2eff83b"; -- 2733635643
        operand2 <= x"348cadd9"; -- 881634777
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4fcd5e41"; -- 1338859073
        operand2 <= x"950ca799"; -- 2500634521
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4fcd5e41"; -- 1338859073
        operand2 <= x"950ca799"; -- 2500634521
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5c77cfdf"; -- 1551355871
        operand2 <= x"36ff231c"; -- 922690332
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5c77cfdf"; -- 1551355871
        operand2 <= x"36ff231c"; -- 922690332
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f1d96c30"; -- 4057558064
        operand2 <= x"fce0ffff"; -- 4242604031
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f1d96c30"; -- 4057558064
        operand2 <= x"fce0ffff"; -- 4242604031
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"42eb057d"; -- 1122698621
        operand2 <= x"0b37886d"; -- 188188781
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"42eb057d"; -- 1122698621
        operand2 <= x"0b37886d"; -- 188188781
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"647ad0a7"; -- 1685770407
        operand2 <= x"0eb1e22e"; -- 246538798
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"647ad0a7"; -- 1685770407
        operand2 <= x"0eb1e22e"; -- 246538798
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"afd5c8ac"; -- 2950023340
        operand2 <= x"c50c9e9f"; -- 3305938591
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"afd5c8ac"; -- 2950023340
        operand2 <= x"c50c9e9f"; -- 3305938591
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5cac8885"; -- 1554811013
        operand2 <= x"e38e7122"; -- 3817763106
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5cac8885"; -- 1554811013
        operand2 <= x"e38e7122"; -- 3817763106
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"34a856f8"; -- 883447544
        operand2 <= x"dc365a78"; -- 3694549624
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"34a856f8"; -- 883447544
        operand2 <= x"dc365a78"; -- 3694549624
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"453337aa"; -- 1160984490
        operand2 <= x"9004b2d6"; -- 2416227030
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"453337aa"; -- 1160984490
        operand2 <= x"9004b2d6"; -- 2416227030
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"760df6c8"; -- 1980626632
        operand2 <= x"701342d8"; -- 1880310488
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"760df6c8"; -- 1980626632
        operand2 <= x"701342d8"; -- 1880310488
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"54ab885e"; -- 1420527710
        operand2 <= x"94a4f181"; -- 2493837697
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"54ab885e"; -- 1420527710
        operand2 <= x"94a4f181"; -- 2493837697
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b4985f88"; -- 3029884808
        operand2 <= x"ca486a8b"; -- 3393743499
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b4985f88"; -- 3029884808
        operand2 <= x"ca486a8b"; -- 3393743499
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fa15952e"; -- 4195718446
        operand2 <= x"6b84c93d"; -- 1803864381
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fa15952e"; -- 4195718446
        operand2 <= x"6b84c93d"; -- 1803864381
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f767964f"; -- 4150761039
        operand2 <= x"b3bfef81"; -- 3015700353
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f767964f"; -- 4150761039
        operand2 <= x"b3bfef81"; -- 3015700353
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1d2f7045"; -- 489648197
        operand2 <= x"a720e998"; -- 2803952024
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1d2f7045"; -- 489648197
        operand2 <= x"a720e998"; -- 2803952024
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1e239a58"; -- 505649752
        operand2 <= x"00f1e1d1"; -- 15851985
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1e239a58"; -- 505649752
        operand2 <= x"00f1e1d1"; -- 15851985
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2bb590dc"; -- 733319388
        operand2 <= x"7ca1c70a"; -- 2090977034
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2bb590dc"; -- 733319388
        operand2 <= x"7ca1c70a"; -- 2090977034
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dd9f7880"; -- 3718215808
        operand2 <= x"b6d664c7"; -- 3067503815
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dd9f7880"; -- 3718215808
        operand2 <= x"b6d664c7"; -- 3067503815
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b07bd762"; -- 2960906082
        operand2 <= x"f673a071"; -- 4134772849
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b07bd762"; -- 2960906082
        operand2 <= x"f673a071"; -- 4134772849
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"25a477df"; -- 631535583
        operand2 <= x"ba7675de"; -- 3128325598
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"25a477df"; -- 631535583
        operand2 <= x"ba7675de"; -- 3128325598
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ba26267f"; -- 3123062399
        operand2 <= x"e2110f59"; -- 3792768857
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ba26267f"; -- 3123062399
        operand2 <= x"e2110f59"; -- 3792768857
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3e421b8c"; -- 1044519820
        operand2 <= x"3a609fb8"; -- 979410872
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3e421b8c"; -- 1044519820
        operand2 <= x"3a609fb8"; -- 979410872
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"db0ec4f6"; -- 3675178230
        operand2 <= x"69b46e50"; -- 1773432400
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"db0ec4f6"; -- 3675178230
        operand2 <= x"69b46e50"; -- 1773432400
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"414292fa"; -- 1094882042
        operand2 <= x"98af6562"; -- 2561631586
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"414292fa"; -- 1094882042
        operand2 <= x"98af6562"; -- 2561631586
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"49201351"; -- 1226838865
        operand2 <= x"52b7904e"; -- 1387761742
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"49201351"; -- 1226838865
        operand2 <= x"52b7904e"; -- 1387761742
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3e0daabf"; -- 1041083071
        operand2 <= x"a82daaf5"; -- 2821565173
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3e0daabf"; -- 1041083071
        operand2 <= x"a82daaf5"; -- 2821565173
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"acd1f95a"; -- 2899442010
        operand2 <= x"01f7dcd8"; -- 33021144
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"acd1f95a"; -- 2899442010
        operand2 <= x"01f7dcd8"; -- 33021144
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"df1ef987"; -- 3743349127
        operand2 <= x"8e785a65"; -- 2390252133
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"df1ef987"; -- 3743349127
        operand2 <= x"8e785a65"; -- 2390252133
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"358fc2b5"; -- 898613941
        operand2 <= x"8be964d7"; -- 2347328727
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"358fc2b5"; -- 898613941
        operand2 <= x"8be964d7"; -- 2347328727
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7b6b68c4"; -- 2070636740
        operand2 <= x"3ce0697b"; -- 1021340027
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7b6b68c4"; -- 2070636740
        operand2 <= x"3ce0697b"; -- 1021340027
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9135e6d1"; -- 2436228817
        operand2 <= x"e373496d"; -- 3815983469
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '1';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9135e6d1"; -- 2436228817
        operand2 <= x"e373496d"; -- 3815983469
        ALUOp <= "011";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f4ab81f5"; -- 4104880629
        operand2 <= x"e96851ef"; -- 3915928047
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"de13d3e4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3e1da5f0"; -- 1042130416
        operand2 <= x"78a0fe1c"; -- 2023816732
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b6bea40c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"449fedf0"; -- 1151331824
        operand2 <= x"3625294a"; -- 908405066
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7ac5173a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"93300a89"; -- 2469399177
        operand2 <= x"15574928"; -- 358041896
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a88753b1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a602dca5"; -- 2785205413
        operand2 <= x"bf0ce31f"; -- 3205292831
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"650fbfc4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"284bdc22"; -- 676060194
        operand2 <= x"2650ac52"; -- 642821202
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4e9c8874" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d977463b"; -- 3648472635
        operand2 <= x"d6b7d8e7"; -- 3602372839
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b02f1f22" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c4734a51"; -- 3295890001
        operand2 <= x"0096227f"; -- 9839231
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c5096cd0" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d9cda202"; -- 3654132226
        operand2 <= x"4c7c3d24"; -- 1283210532
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2649df26" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8ecc5f2e"; -- 2395758382
        operand2 <= x"477650c3"; -- 1198936259
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d642aff1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fd1b5b04"; -- 4246428420
        operand2 <= x"b3a58f69"; -- 3013971817
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b0c0ea6d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4af7b5e9"; -- 1257747945
        operand2 <= x"bed4f6d5"; -- 3201627861
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"09ccacbe" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2e3a7c16"; -- 775584790
        operand2 <= x"34096deb"; -- 873033195
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6243ea01" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e424918b"; -- 3827601803
        operand2 <= x"b1094943"; -- 2970175811
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"952ddace" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"96d70a67"; -- 2530675303
        operand2 <= x"480e0e3b"; -- 1208880699
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"dee518a2" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6607b86e"; -- 1711781998
        operand2 <= x"a024900e"; -- 2686750734
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"062c487c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"646b3396"; -- 1684747158
        operand2 <= x"22fd9a43"; -- 587045443
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8768cdd9" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c38e53dc"; -- 3280884700
        operand2 <= x"13314680"; -- 321996416
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d6bf9a5c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4d5af1ca"; -- 1297805770
        operand2 <= x"5810821d"; -- 1477476893
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a56b73e7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"362b22cd"; -- 908796621
        operand2 <= x"21fd1c8e"; -- 570236046
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"58283f5b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7ba9c771"; -- 2074724209
        operand2 <= x"fcb00737"; -- 4239394615
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7859cea8" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"be4ece17"; -- 3192835607
        operand2 <= x"fe313d24"; -- 4264639780
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bc800b3b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"78608d61"; -- 2019593569
        operand2 <= x"16c3a418"; -- 381920280
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8f243179" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"daf6885f"; -- 3673589855
        operand2 <= x"cd308b1a"; -- 3442510618
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a8271379" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2a001d3f"; -- 704650559
        operand2 <= x"89079658"; -- 2298975832
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b307b397" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6d62b227"; -- 1835184679
        operand2 <= x"228e8c30"; -- 579767344
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8ff13e57" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7532cb61"; -- 1966263137
        operand2 <= x"ad764f89"; -- 2910211977
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"22a91aea" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f943dfa9"; -- 4181974953
        operand2 <= x"53a772ac"; -- 1403482796
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4ceb5255" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e6a093fc"; -- 3869283324
        operand2 <= x"df19463d"; -- 3742975549
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c5b9da39" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"407341e5"; -- 1081295333
        operand2 <= x"925274cc"; -- 2454877388
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d2c5b6b1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1404dcc3"; -- 335862979
        operand2 <= x"74fa07ec"; -- 1962543084
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"88fee4af" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"36ec3541"; -- 921449793
        operand2 <= x"9a1a17e3"; -- 2585401315
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d1064d24" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9aaca1d8"; -- 2595004888
        operand2 <= x"ce1f6807"; -- 3458164743
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"68cc09df" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4d03faaf"; -- 1292106415
        operand2 <= x"68b0c378"; -- 1756414840
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b5b4be27" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9343ec59"; -- 2470702169
        operand2 <= x"71777144"; -- 1903653188
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"04bb5d9d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"12194591"; -- 303646097
        operand2 <= x"e7e1abb3"; -- 3890326451
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f9faf144" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7e36c6f3"; -- 2117519091
        operand2 <= x"9a59fd91"; -- 2589588881
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1890c484" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dae325fc"; -- 3672319484
        operand2 <= x"63bc70cb"; -- 1673294027
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3e9f96c7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d0512a6c"; -- 3494980204
        operand2 <= x"ae01c86d"; -- 2919352429
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7e52f2d9" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5ddace10"; -- 1574620688
        operand2 <= x"40faaad6"; -- 1090169558
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9ed578e6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3e21de82"; -- 1042407042
        operand2 <= x"f2c0d2bf"; -- 4072723135
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"30e2b141" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4180adca"; -- 1098952138
        operand2 <= x"6201ae30"; -- 1644277296
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a3825bfa" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bf5b7df9"; -- 3210444281
        operand2 <= x"ffd7a52d"; -- 4292322605
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bf332326" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1c521f1e"; -- 475143966
        operand2 <= x"20a34977"; -- 547572087
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3cf56895" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d1bb267a"; -- 3518703226
        operand2 <= x"fa16ddf2"; -- 4195802610
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"cbd2046c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a1261c12"; -- 2703629330
        operand2 <= x"74e5d450"; -- 1961219152
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"160bf062" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"151a9617"; -- 354063895
        operand2 <= x"30c361d2"; -- 818110930
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"45ddf7e9" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"aa5e38e5"; -- 2858301669
        operand2 <= x"a6fbe690"; -- 2801526416
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"515a1f75" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"00e30548"; -- 14878024
        operand2 <= x"f7131bcc"; -- 4145224652
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f7f62114" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1c2ddd79"; -- 472767865
        operand2 <= x"6246ae7b"; -- 1648799355
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7e748bf4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ebea1293"; -- 3957985939
        operand2 <= x"6ce1f871"; -- 1826748529
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"58cc0b04" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"836e0a90"; -- 2205026960
        operand2 <= x"5e97243e"; -- 1586963518
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"e2052ece" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"34242206"; -- 874783238
        operand2 <= x"36b76ecc"; -- 917991116
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6adb90d2" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b00bb42d"; -- 2953557037
        operand2 <= x"3f62baf5"; -- 1063434997
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ef6e6f22" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f1587369"; -- 4049105769
        operand2 <= x"b9c3aa21"; -- 3116608033
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ab1c1d8a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1d875727"; -- 495408935
        operand2 <= x"1488a4af"; -- 344499375
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"320ffbd6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"31d04dce"; -- 835734990
        operand2 <= x"8e6d6b6d"; -- 2389535597
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c03db93b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"efda0d89"; -- 4024044937
        operand2 <= x"4ec5ae41"; -- 1321578049
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3e9fbbca" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"908a85cd"; -- 2424997325
        operand2 <= x"0e00b799"; -- 234928025
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9e8b3d66" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ca5cd8d2"; -- 3395082450
        operand2 <= x"cb0810cb"; -- 3406303435
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9564e99d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a8e22fb9"; -- 2833395641
        operand2 <= x"7548738a"; -- 1967682442
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1e2aa343" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"346c1e36"; -- 879500854
        operand2 <= x"6e954ccb"; -- 1855278283
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a3016b01" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"508a6a0f"; -- 1351248399
        operand2 <= x"1e4fbb50"; -- 508541776
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6eda255f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"325e7c76"; -- 845053046
        operand2 <= x"09510b23"; -- 156306211
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3baf8799" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"cde938ae"; -- 3454613678
        operand2 <= x"5132242c"; -- 1362240556
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1f1b5cda" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1bcff4d7"; -- 466613463
        operand2 <= x"883ce303"; -- 2285691651
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a40cd7da" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"97167f11"; -- 2534833937
        operand2 <= x"762a8fef"; -- 1982500847
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0d410f00" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3307ecb2"; -- 856157362
        operand2 <= x"dc7e1069"; -- 3699249257
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0f85fd1b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6594d6bd"; -- 1704253117
        operand2 <= x"285fd2a5"; -- 677368485
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8df4a962" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0705bcf9"; -- 117816569
        operand2 <= x"72cd5b09"; -- 1926060809
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"79d31802" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0aad666b"; -- 179136107
        operand2 <= x"95b54fcc"; -- 2511687628
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a062b637" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"93d19401"; -- 2479985665
        operand2 <= x"0cf04bd6"; -- 217074646
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a0c1dfd7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"13ae0f61"; -- 330174305
        operand2 <= x"da875195"; -- 3666301333
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ee3560f6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"24f132c4"; -- 619786948
        operand2 <= x"a26feb6d"; -- 2725243757
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c7611e31" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7ff066ad"; -- 2146461357
        operand2 <= x"cbd928e3"; -- 3420006627
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4bc98f90" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"18dccf5e"; -- 417124190
        operand2 <= x"997e6ff0"; -- 2575200240
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b25b3f4e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e9ab4b44"; -- 3920317252
        operand2 <= x"a2975cfb"; -- 2727828731
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8c42a83f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"067926d5"; -- 108603093
        operand2 <= x"8ab8b272"; -- 2327360114
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9131d947" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c51da0b5"; -- 3307053237
        operand2 <= x"4e085285"; -- 1309168261
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1325f33a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"49dd3cef"; -- 1239235823
        operand2 <= x"a908f6ee"; -- 2835937006
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f2e633dd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dcb5fd77"; -- 3702914423
        operand2 <= x"6efd3fa3"; -- 1862090659
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4bb33d1a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6d3c548a"; -- 1832670346
        operand2 <= x"a905c2c5"; -- 2835727045
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1642174f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"cc7ee704"; -- 3430868740
        operand2 <= x"c640a8ea"; -- 3326126314
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"92bf8fee" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bc7c5346"; -- 3162264390
        operand2 <= x"3a6a25eb"; -- 980035051
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f6e67931" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d3ab114d"; -- 3551203661
        operand2 <= x"a7de8cf9"; -- 2816380153
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7b899e46" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4adc68f7"; -- 1255958775
        operand2 <= x"864e8dcf"; -- 2253295055
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d12af6c6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f4ab8600"; -- 4104881664
        operand2 <= x"b07ba1ce"; -- 2960892366
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a52727ce" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"63fc5323"; -- 1677480739
        operand2 <= x"f9b06969"; -- 4189088105
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"5dacbc8c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b7688b92"; -- 3077082002
        operand2 <= x"5da14bac"; -- 1570851756
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1509d73e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c516509d"; -- 3306573981
        operand2 <= x"feefe125"; -- 4277133605
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c40631c2" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d1a8ea1b"; -- 3517508123
        operand2 <= x"5da4f865"; -- 1571092581
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2f4de280" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f8c6bebe"; -- 4173774526
        operand2 <= x"e457dc1f"; -- 3830963231
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"dd1e9add" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0f865ab0"; -- 260463280
        operand2 <= x"11a592b5"; -- 296063669
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"212bed65" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5f02bac0"; -- 1594014400
        operand2 <= x"a4503319"; -- 2756719385
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0352edd9" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"09768352"; -- 158761810
        operand2 <= x"51877b3b"; -- 1367833403
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"5afdfe8d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"041ff138"; -- 69202232
        operand2 <= x"ce415d41"; -- 3460390209
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d2614e79" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8f0526d2"; -- 2399479506
        operand2 <= x"a692ec43"; -- 2794646595
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"35981315" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"92ba06c5"; -- 2461664965
        operand2 <= x"20736abb"; -- 544434875
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b32d7180" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8b8d1162"; -- 2341278050
        operand2 <= x"384ed8b0"; -- 944691376
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c3dbea12" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6c51507a"; -- 1817268346
        operand2 <= x"e4ddd78f"; -- 3839743887
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"512f2809" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d5a16c52"; -- 3584126034
        operand2 <= x"bf230bad"; -- 3206745005
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"94c477ff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"325561b1"; -- 844456369
        operand2 <= x"0b5418a3"; -- 190060707
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3da97a54" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fbb9b329"; -- 4223251241
        operand2 <= x"0ca182a0"; -- 211911328
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"085b35c9" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f5c17254"; -- 4123095636
        operand2 <= x"1a6288ec"; -- 442665196
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1023fb40" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0989df91"; -- 160030609
        operand2 <= x"fe320b45"; -- 4264692549
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"07bbead6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"cc0b50c1"; -- 3423293633
        operand2 <= x"bb66ff07"; -- 3144089351
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"87724fc8" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a1eee493"; -- 2716787859
        operand2 <= x"bca03567"; -- 3164616039
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"5e8f19fa" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"256fa88f"; -- 628074639
        operand2 <= x"8e026a93"; -- 2382523027
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b3721322" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c3e41a74"; -- 3286506100
        operand2 <= x"8e676c42"; -- 2389142594
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"524b86b6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5e0d8b46"; -- 1577945926
        operand2 <= x"65b4c119"; -- 1706344729
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c3c24c5f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2a349f3a"; -- 708091706
        operand2 <= x"9694f31f"; -- 2526343967
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c0c99259" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9c463165"; -- 2621845861
        operand2 <= x"b0b81f7c"; -- 2964856700
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4cfe50e1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1d5f5801"; -- 492787713
        operand2 <= x"94825475"; -- 2491569269
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b1e1ac76" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7f829064"; -- 2139263076
        operand2 <= x"4a14ce31"; -- 1242877489
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c9975e95" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e71a1976"; -- 3877247350
        operand2 <= x"38d9c75b"; -- 953796443
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1ff3e0d1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"77a8f766"; -- 2007562086
        operand2 <= x"0fde4de1"; -- 266227169
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"87874547" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"01edb1ab"; -- 32354731
        operand2 <= x"f708667e"; -- 4144522878
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f8f61829" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2aff6b62"; -- 721382242
        operand2 <= x"f1d966aa"; -- 4057556650
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1cd8d20c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2b41c2cd"; -- 725729997
        operand2 <= x"23cf5ea3"; -- 600792739
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4f112170" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"abf3f4c0"; -- 2884891840
        operand2 <= x"e934242b"; -- 3912508459
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"952818eb" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c65252b7"; -- 3327283895
        operand2 <= x"f678da34"; -- 4135115316
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bccb2ceb" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"71db2f4b"; -- 1910189899
        operand2 <= x"cd887c12"; -- 3448273938
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3f63ab5d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3d9ca30c"; -- 1033675532
        operand2 <= x"e825d9f4"; -- 3894794740
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"25c27d00" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"cb4cd967"; -- 3410811239
        operand2 <= x"b3bc915c"; -- 3015479644
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7f096ac3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1de64d39"; -- 501632313
        operand2 <= x"4c921141"; -- 1284641089
        ALUOp <= "100";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6a785e7a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"526c8b64"; -- 1382845284
        operand2 <= x"dd8003d7"; -- 3716154327
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"74ec878d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dcc0c228"; -- 3703620136
        operand2 <= x"e0a21441"; -- 3768718401
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fc1eade7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"96c49e12"; -- 2529467922
        operand2 <= x"83adf42b"; -- 2209215531
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1316a9e7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"45bc9b54"; -- 1169988436
        operand2 <= x"7487f8e6"; -- 1955068134
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d134a26e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2c484640"; -- 742934080
        operand2 <= x"08b0f977"; -- 145815927
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"23974cc9" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ab5cf1b8"; -- 2874995128
        operand2 <= x"d5eea07c"; -- 3589185660
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d56e513c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"aefddb99"; -- 2935872409
        operand2 <= x"713f9c74"; -- 1899994228
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3dbe3f25" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a430e71e"; -- 2754668318
        operand2 <= x"07ece2d2"; -- 132965074
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9c44044c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"acd60a65"; -- 2899708517
        operand2 <= x"5fa71f91"; -- 1604788113
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4d2eead4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"76a62804"; -- 1990600708
        operand2 <= x"2321896b"; -- 589400427
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"53849e99" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1d1cdea3"; -- 488431267
        operand2 <= x"f3d9f157"; -- 4091146583
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2942ed4c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"10450dfe"; -- 272961022
        operand2 <= x"f76e222b"; -- 4151190059
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"18d6ebd3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9f628924"; -- 2674034980
        operand2 <= x"98943442"; -- 2559849538
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"06ce54e2" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"956db9d1"; -- 2506996177
        operand2 <= x"794bdfba"; -- 2035015610
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1c21da17" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b029d724"; -- 2955532068
        operand2 <= x"fe09bb7e"; -- 4262050686
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b2201ba6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9fc73c9f"; -- 2680634527
        operand2 <= x"41b68ee1"; -- 1102483169
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"5e10adbe" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2a535c59"; -- 710106201
        operand2 <= x"2b7c3392"; -- 729559954
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fed728c7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bb426949"; -- 3141691721
        operand2 <= x"ead2f1b7"; -- 3939692983
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d06f7792" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1fa8f64a"; -- 531166794
        operand2 <= x"2f5008c0"; -- 793774272
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f058ed8a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a004b0ff"; -- 2684662015
        operand2 <= x"b1428295"; -- 2973926037
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"eec22e6a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"781a615b"; -- 2014994779
        operand2 <= x"85fc9662"; -- 2247923298
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f21dcaf9" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a3ce8c10"; -- 2748222480
        operand2 <= x"b1c152fa"; -- 2982236922
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f20d3916" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"20d59718"; -- 550868760
        operand2 <= x"a39d099b"; -- 2744977819
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7d388d7d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f1d101b3"; -- 4057006515
        operand2 <= x"6b6af8e4"; -- 1802172644
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"866608cf" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"269720d1"; -- 647438545
        operand2 <= x"e8ea5d97"; -- 3907673495
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3dacc33a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3753d2ba"; -- 928240314
        operand2 <= x"feeb93fb"; -- 4276851707
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"38683ebf" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a81d44fc"; -- 2820490492
        operand2 <= x"c6bbe971"; -- 3334203761
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"e1615b8b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4c0b6bed"; -- 1275816941
        operand2 <= x"6e0b503d"; -- 1846235197
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"de001bb0" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0195436a"; -- 26559338
        operand2 <= x"c5874d98"; -- 3313978776
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3c0df5d2" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8209caae"; -- 2181679790
        operand2 <= x"3021ca2d"; -- 807520813
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"51e80081" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fe5afe5f"; -- 4267376223
        operand2 <= x"b3744cb5"; -- 3010743477
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4ae6b1aa" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3dfbb049"; -- 1039904841
        operand2 <= x"e3fa7944"; -- 3824843076
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"5a013705" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5bea9f19"; -- 1542102809
        operand2 <= x"928ddae7"; -- 2458770151
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c95cc432" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"968decfe"; -- 2525883646
        operand2 <= x"fbe4257d"; -- 4226033021
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9aa9c781" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"eb3a7af7"; -- 3946478327
        operand2 <= x"1b62f1ad"; -- 459469229
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"cfd7894a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"01b07d49"; -- 28343625
        operand2 <= x"28bbbd54"; -- 683392340
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d8f4bff5" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c25e0916"; -- 3260942614
        operand2 <= x"2a552bed"; -- 710224877
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9808dd29" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5eaf2cf4"; -- 1588538612
        operand2 <= x"a392ce71"; -- 2744307313
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"bb1c5e83" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"242c9382"; -- 606901122
        operand2 <= x"48180366"; -- 1209533286
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"dc14901c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"71ebc56f"; -- 1911276911
        operand2 <= x"f8ab355e"; -- 4171969886
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"79409011" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a21aa3a3"; -- 2719654819
        operand2 <= x"5fa94342"; -- 1604928322
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"42716061" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"67690d4b"; -- 1734937931
        operand2 <= x"d7900513"; -- 3616539923
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8fd90838" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3a5f1edc"; -- 979312348
        operand2 <= x"00ff2ad7"; -- 16722647
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"395ff405" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8a95da25"; -- 2325076517
        operand2 <= x"e5a22ccf"; -- 3852610767
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a4f3ad56" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"646a2b12"; -- 1684679442
        operand2 <= x"01ad7a32"; -- 28146226
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"62bcb0e0" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4e8318ab"; -- 1317214379
        operand2 <= x"fa3d28bd"; -- 4198312125
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"5445efee" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e75cab3d"; -- 3881610045
        operand2 <= x"adeb113c"; -- 2917863740
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"39719a01" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"80f5671f"; -- 2163566367
        operand2 <= x"4f475f6d"; -- 1330077549
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"31ae07b2" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9042ae93"; -- 2420289171
        operand2 <= x"8ce0949b"; -- 2363528347
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"036219f8" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8dd24781"; -- 2379368321
        operand2 <= x"3ab4bf71"; -- 984924017
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"531d8810" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"62160fa2"; -- 1645612962
        operand2 <= x"59f6ac1c"; -- 1509338140
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"081f6386" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"120608c1"; -- 302385345
        operand2 <= x"5118450d"; -- 1360545037
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c0edc3b4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8af9a6a8"; -- 2331616936
        operand2 <= x"07cd383f"; -- 130889791
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"832c6e69" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b2361c9d"; -- 2989890717
        operand2 <= x"db0be549"; -- 3674989897
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d72a3754" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"47dadc14"; -- 1205525524
        operand2 <= x"ea8a5982"; -- 3934935426
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"5d508292" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1d1d8a1e"; -- 488475166
        operand2 <= x"6516b49f"; -- 1695986847
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b806d57f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"87dd36ac"; -- 2279421612
        operand2 <= x"da408800"; -- 3661662208
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ad9caeac" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1d5b9e90"; -- 492543632
        operand2 <= x"9746b7aa"; -- 2537994154
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8614e6e6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f7a48334"; -- 4154753844
        operand2 <= x"f16bd5c9"; -- 4050376137
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0638ad6b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"24f33063"; -- 619917411
        operand2 <= x"251cc623"; -- 622642723
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffd66a40" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"95766b4d"; -- 2507565901
        operand2 <= x"da88cdff"; -- 3666398719
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"baed9d4e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3540068a"; -- 893388426
        operand2 <= x"1a1dd734"; -- 438163252
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1b222f56" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"18e8d3fd"; -- 417911805
        operand2 <= x"e8394977"; -- 3896068471
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"30af8a86" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7ddc1075"; -- 2111574133
        operand2 <= x"5d2c5169"; -- 1563185513
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"20afbf0c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ea41c45e"; -- 3930178654
        operand2 <= x"bea52ab2"; -- 3198495410
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2b9c99ac" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"65ebda42"; -- 1709955650
        operand2 <= x"cc221131"; -- 3424784689
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"99c9c911" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"48b02ed0"; -- 1219505872
        operand2 <= x"39d557e2"; -- 970282978
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0edad6ee" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"41f1e060"; -- 1106370656
        operand2 <= x"156d53a9"; -- 359486377
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2c848cb7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d4e2eb94"; -- 3571641236
        operand2 <= x"6a62bb5c"; -- 1784855388
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6a803038" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e05611cb"; -- 3763737035
        operand2 <= x"ec0f9a69"; -- 3960445545
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f4467762" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1ffcd708"; -- 536663816
        operand2 <= x"04912401"; -- 76620801
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1b6bb307" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"de85e77a"; -- 3733317498
        operand2 <= x"d19b7b75"; -- 3516627829
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0cea6c05" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d600d5d9"; -- 3590378969
        operand2 <= x"89604ada"; -- 2304789210
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4ca08aff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d42c8762"; -- 3559688034
        operand2 <= x"5f6b5573"; -- 1600869747
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"74c131ef" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0f413b38"; -- 255933240
        operand2 <= x"6cba2d5a"; -- 1824140634
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a2870dde" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7391ce01"; -- 1938935297
        operand2 <= x"8f399499"; -- 2402915481
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"e4583968" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d50fb07e"; -- 3574575230
        operand2 <= x"5d4ef244"; -- 1565454916
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"77c0be3a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"66964746"; -- 1721124678
        operand2 <= x"6d7c9723"; -- 1836881699
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f919b023" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"94812847"; -- 2491492423
        operand2 <= x"9c4e9262"; -- 2622394978
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f83295e5" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"39179fed"; -- 957849581
        operand2 <= x"8a7f8c02"; -- 2323614722
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ae9813eb" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"597155a5"; -- 1500599717
        operand2 <= x"143cd0f9"; -- 339529977
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"453484ac" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"615e01cb"; -- 1633550795
        operand2 <= x"3095c4ce"; -- 815121614
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"30c83cfd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4b7b1aea"; -- 1266359018
        operand2 <= x"6cbce155"; -- 1824317781
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"debe3995" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"128daae3"; -- 311274211
        operand2 <= x"0ff1e1d6"; -- 267510230
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"029bc90d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0ebb14c0"; -- 247141568
        operand2 <= x"0a3e1fa0"; -- 171843488
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"047cf520" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2be56df1"; -- 736456177
        operand2 <= x"6d82bfa8"; -- 1837285288
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"be62ae49" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"443d8560"; -- 1144882528
        operand2 <= x"a99d839f"; -- 2845672351
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9aa001c1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f8301caa"; -- 4163902634
        operand2 <= x"4e6dd277"; -- 1315820151
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a9c24a33" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"83859f9a"; -- 2206572442
        operand2 <= x"44edbe4d"; -- 1156431437
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3e97e14d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0e0691f7"; -- 235311607
        operand2 <= x"a252a464"; -- 2723325028
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6bb3ed93" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c72f7f3d"; -- 3341778749
        operand2 <= x"f5dc6e99"; -- 4124864153
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d15310a4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e9d187ae"; -- 3922823086
        operand2 <= x"b149875c"; -- 2974386012
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"38880052" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d745a34c"; -- 3611665228
        operand2 <= x"33906859"; -- 865101913
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a3b53af3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f3c387e6"; -- 4089677798
        operand2 <= x"a54f9b20"; -- 2773457696
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4e73ecc6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fa1c8f9f"; -- 4196175775
        operand2 <= x"64eeae46"; -- 1693363782
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"952de159" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0b0b031d"; -- 185271069
        operand2 <= x"612f223b"; -- 1630478907
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a9dbe0e2" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f51fba67"; -- 4112497255
        operand2 <= x"97c4d12a"; -- 2546258218
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"5d5ae93d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e2ba63a1"; -- 3803866017
        operand2 <= x"bd636083"; -- 3177406595
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2557031e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a94ec78b"; -- 2840512395
        operand2 <= x"cb344723"; -- 3409200931
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"de1a8068" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7bee9327"; -- 2079232807
        operand2 <= x"37b3a6c0"; -- 934520512
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"443aec67" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"73f83b20"; -- 1945647904
        operand2 <= x"e8e7ec64"; -- 3907513444
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8b104ebc" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1bd435ef"; -- 466892271
        operand2 <= x"b976e69d"; -- 3111577245
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"625d4f52" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8109e721"; -- 2164909857
        operand2 <= x"05f96e5a"; -- 100232794
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7b1078c7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"500be60d"; -- 1342957069
        operand2 <= x"744d1a88"; -- 1951210120
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"dbbecb85" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"85582247"; -- 2237145671
        operand2 <= x"fb95567a"; -- 4220868218
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"89c2cbcd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f670b834"; -- 4134582324
        operand2 <= x"d9825621"; -- 3649197601
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1cee6213" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"990611b9"; -- 2567311801
        operand2 <= x"ca3f461f"; -- 3393144351
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"cec6cb9a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"452b3995"; -- 1160460693
        operand2 <= x"28b31e19"; -- 682827289
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1c781b7c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7b383e58"; -- 2067283544
        operand2 <= x"eda972bc"; -- 3987305148
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8d8ecb9c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fa36cc33"; -- 4197895219
        operand2 <= x"11013f79"; -- 285294457
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"e9358cba" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"427fe395"; -- 1115677589
        operand2 <= x"fe83e838"; -- 4270057528
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"43fbfb5d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"78f475c5"; -- 2029286853
        operand2 <= x"75e158ad"; -- 1977702573
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"03131d18" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8db4017d"; -- 2377384317
        operand2 <= x"c0217a63"; -- 3223419491
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"cd92871a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9928db21"; -- 2569591585
        operand2 <= x"2581f1d7"; -- 629273047
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"73a6e94a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"be7c0ca8"; -- 3195800744
        operand2 <= x"4c899bcd"; -- 1284086733
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"71f270db" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a4ec932c"; -- 2766967596
        operand2 <= x"ab459b43"; -- 2873465667
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f9a6f7e9" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a4765560"; -- 2759218528
        operand2 <= x"0a7f617b"; -- 176120187
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"99f6f3e5" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"92691ffd"; -- 2456363005
        operand2 <= x"51ebed2a"; -- 1374416170
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"407d32d3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"78f83428"; -- 2029532200
        operand2 <= x"f16c1535"; -- 4050392373
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"878c1ef3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1fba9020"; -- 532320288
        operand2 <= x"36e38b07"; -- 920881927
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"e8d70519" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1c44b06b"; -- 474263659
        operand2 <= x"f5bba5ff"; -- 4122715647
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"26890a6c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6993441c"; -- 1771258908
        operand2 <= x"01bc3e91"; -- 29114001
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"67d7058b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6c0d7d81"; -- 1812823425
        operand2 <= x"794b04ea"; -- 2034959594
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f2c27897" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d0979af8"; -- 3499596536
        operand2 <= x"3102cbb9"; -- 822266809
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9f94cf3f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2ad3de2f"; -- 718528047
        operand2 <= x"46e6f502"; -- 1189541122
        ALUOp <= "101";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"e3ece92d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0c9060a9"; -- 210788521
        operand2 <= x"83736247"; -- 2205377095
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"48305480" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"43ac1119"; -- 1135350041
        operand2 <= x"c3962fed"; -- 3281399789
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"82232000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"425ab61a"; -- 1113241114
        operand2 <= x"c33614b9"; -- 3275101369
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"34000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b23f9ecc"; -- 2990513868
        operand2 <= x"f4ab72fc"; -- 4104876796
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c0000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"47ad927a"; -- 1202557562
        operand2 <= x"7a1ca299"; -- 2048696985
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f4000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2565e40d"; -- 627434509
        operand2 <= x"a3f41263"; -- 2750681699
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2b2f2068" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"45ea7231"; -- 1172992561
        operand2 <= x"3f5a6df2"; -- 1062890994
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c8c40000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4eab32c1"; -- 1319842497
        operand2 <= x"a12e563a"; -- 2704168506
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"04000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a50ffac3"; -- 2769287875
        operand2 <= x"cf51cbdd"; -- 3478244317
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"60000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2cf438aa"; -- 754202794
        operand2 <= x"0ac2f8b4"; -- 180549812
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8aa00000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9b4aefe6"; -- 2605379558
        operand2 <= x"06dc2357"; -- 115090263
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f3000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"19536d01"; -- 424897793
        operand2 <= x"f54fb9bc"; -- 4115642812
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"10000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e98a0104"; -- 3918135556
        operand2 <= x"8d770b3a"; -- 2373389114
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"10000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"89fd3d73"; -- 2315074931
        operand2 <= x"54b2491d"; -- 1420970269
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"60000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ebbe1464"; -- 3955102820
        operand2 <= x"ef1a0efa"; -- 4011462394
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"90000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4aecb921"; -- 1257027873
        operand2 <= x"c3261283"; -- 3274052227
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"5765c908" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"86ba2099"; -- 2260344985
        operand2 <= x"40a0f26a"; -- 1084289642
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"e8826400" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9fb4a81c"; -- 2679416860
        operand2 <= x"3625f464"; -- 908457060
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fb4a81c0" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"46d92937"; -- 1188636983
        operand2 <= x"3f1f49e4"; -- 1059015140
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6d929370" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0cd11c4b"; -- 215030859
        operand2 <= x"95faf554"; -- 2516251988
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c4b00000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9c80f34c"; -- 2625696588
        operand2 <= x"02b95a04"; -- 45701636
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c80f34c0" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"65716655"; -- 1701930581
        operand2 <= x"29a55bce"; -- 698702798
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"59954000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d3b197c5"; -- 3551631301
        operand2 <= x"6fe7bec8"; -- 1877458632
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b197c500" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8a2e7e28"; -- 2318302760
        operand2 <= x"46eb9064"; -- 1189843044
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a2e7e280" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9971b9dc"; -- 2574367196
        operand2 <= x"a56dc373"; -- 2775434099
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"cee00000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"26ede8f2"; -- 653125874
        operand2 <= x"adb52007"; -- 2914328583
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"76f47900" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dd0d1a01"; -- 3708623361
        operand2 <= x"bad0d05b"; -- 3134247003
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"08000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"893ce086"; -- 2302468230
        operand2 <= x"218d4568"; -- 562906472
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3ce08600" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6ec0ef30"; -- 1858137904
        operand2 <= x"a529200e"; -- 2770935822
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3bcc0000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4258791a"; -- 1113094426
        operand2 <= x"2396d434"; -- 597087284
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"91a00000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"61159106"; -- 1628803334
        operand2 <= x"95482a09"; -- 2504534537
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2b220c00" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e8b2b060"; -- 3904024672
        operand2 <= x"c4f3c014"; -- 3304308756
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"06000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"363f87b9"; -- 910133177
        operand2 <= x"2e485570"; -- 776492400
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"87b90000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"591bc8f5"; -- 1494993141
        operand2 <= x"fd883a03"; -- 4253563395
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c8de47a8" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ed3cc02d"; -- 3980181549
        operand2 <= x"67ffa389"; -- 1744806793
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"79805a00" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fc6c4055"; -- 4234952789
        operand2 <= x"313bce80"; -- 826003072
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fc6c4055" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5cde7965"; -- 1558083941
        operand2 <= x"89478e85"; -- 2303168133
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9bcf2ca0" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6d0a0d08"; -- 1829375240
        operand2 <= x"fce002a4"; -- 4242539172
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d0a0d080" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e020c22e"; -- 3760243246
        operand2 <= x"28e162a5"; -- 685859493
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"041845c0" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"08b1e6e6"; -- 145876710
        operand2 <= x"9e62aebd"; -- 2657267389
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c0000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a1b6e348"; -- 2713117512
        operand2 <= x"b794ef00"; -- 3079991040
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a1b6e348" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3708a313"; -- 923312915
        operand2 <= x"9984d3ef"; -- 2575619055
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"51898000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c2be3e21"; -- 3267247649
        operand2 <= x"3b0d8b7d"; -- 990743421
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"20000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"49dab8f1"; -- 1239070961
        operand2 <= x"76eef5e0"; -- 1995372000
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"49dab8f1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"803835e3"; -- 2151167459
        operand2 <= x"759bf03a"; -- 1973153850
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8c000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"17eccf43"; -- 401395523
        operand2 <= x"ebdc19d9"; -- 3957070297
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"86000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9eb0c928"; -- 2662385960
        operand2 <= x"20405795"; -- 541087637
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"25000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"24ded17c"; -- 618582396
        operand2 <= x"5c500531"; -- 1548748081
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a2f80000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"12a1b3f5"; -- 312587253
        operand2 <= x"edfcd5d1"; -- 3992770001
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"67ea0000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c93a5ea5"; -- 3376045733
        operand2 <= x"2df5127c"; -- 771035772
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"50000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"93737d47"; -- 2473819463
        operand2 <= x"d90cda7f"; -- 3641498239
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"80000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6c14a6d2"; -- 1813292754
        operand2 <= x"8deff63e"; -- 2381313598
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"80000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0aab9151"; -- 179016017
        operand2 <= x"a0f457e0"; -- 2700367840
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0aab9151" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2eedccb7"; -- 787336375
        operand2 <= x"c6929b49"; -- 3331496777
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"db996e00" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"806a068e"; -- 2154432142
        operand2 <= x"b5aba013"; -- 3047923731
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"34700000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8b46a1f7"; -- 2336662007
        operand2 <= x"b0da43b4"; -- 2967094196
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1f700000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"25b17728"; -- 632387368
        operand2 <= x"b564d60b"; -- 3043284491
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"8bb94000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"be0a6954"; -- 3188353364
        operand2 <= x"abfca148"; -- 2885460296
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0a695400" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5b45d786"; -- 1531303814
        operand2 <= x"adfc69e3"; -- 2919000547
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"da2ebc30" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"84648e6a"; -- 2221182570
        operand2 <= x"167abe83"; -- 377142915
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"23247350" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0fa34f1a"; -- 262360858
        operand2 <= x"a208d9dc"; -- 2718489052
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a0000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7cfa566d"; -- 2096780909
        operand2 <= x"c2219c07"; -- 3256982535
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7d2b3680" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d4e00f0b"; -- 3571453707
        operand2 <= x"5238c49d"; -- 1379452061
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"60000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8cd7685b"; -- 2362927195
        operand2 <= x"2d96e762"; -- 764864354
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"335da16c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"854314a6"; -- 2235765926
        operand2 <= x"1984a53e"; -- 428123454
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"80000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"64f5b21d"; -- 1693823517
        operand2 <= x"b3a1b490"; -- 3013719184
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b21d0000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bbfdf1ed"; -- 3153981933
        operand2 <= x"7a872197"; -- 2055676311
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f6800000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6f3f8ddd"; -- 1866436061
        operand2 <= x"eee2deea"; -- 4007845610
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fe377400" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ee49e663"; -- 3997820515
        operand2 <= x"a7547383"; -- 2807329667
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"724f3318" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d2b3e4f7"; -- 3535004919
        operand2 <= x"9484cac5"; -- 2491730629
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"567c9ee0" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"37622ba7"; -- 929180583
        operand2 <= x"932a17f0"; -- 2469009392
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2ba70000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"174d4fef"; -- 390942703
        operand2 <= x"3ad00255"; -- 986710613
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fde00000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"11ac82c8"; -- 296518344
        operand2 <= x"a6fa6d33"; -- 2801429811
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"16400000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bd6e06c4"; -- 3178104516
        operand2 <= x"2dcbe6ff"; -- 768337663
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"36b60151"; -- 917897553
        operand2 <= x"2e75eb33"; -- 779479859
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0a880000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f5869310"; -- 4119237392
        operand2 <= x"ab3a3e48"; -- 2872720968
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"86931000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"957333e5"; -- 2507355109
        operand2 <= x"064f37df"; -- 105854943
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"80000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9a8cf416"; -- 2592928790
        operand2 <= x"881fd17e"; -- 2283786622
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"80000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fb314642"; -- 4214310466
        operand2 <= x"e6b2fe4c"; -- 3870490188
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"14642000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e15ddb9f"; -- 3781024671
        operand2 <= x"d6f1dc28"; -- 3606174760
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"5ddb9f00" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e2e228b3"; -- 3806472371
        operand2 <= x"af8b5b1c"; -- 2945145628
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"30000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"10dd23fb"; -- 282928123
        operand2 <= x"d2d6f2e7"; -- 3537302247
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6e91fd80" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9741af6e"; -- 2537664366
        operand2 <= x"1eb2a776"; -- 515024758
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"db800000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3251c7f4"; -- 844220404
        operand2 <= x"480f2620"; -- 1208952352
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3251c7f4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"41de92d3"; -- 1105105619
        operand2 <= x"a6211c10"; -- 2787187728
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"92d30000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8ea44b90"; -- 2393131920
        operand2 <= x"04d71c25"; -- 81206309
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d4897200" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0fcb672c"; -- 264988460
        operand2 <= x"519f0589"; -- 1369376137
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"96ce5800" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0bb7318a"; -- 196555146
        operand2 <= x"6e490151"; -- 1850278225
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"63140000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b2a580ef"; -- 2997190895
        operand2 <= x"44524f3f"; -- 1146244927
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"80000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6a229bfe"; -- 1780653054
        operand2 <= x"953c8336"; -- 2503770934
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ff800000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3386201c"; -- 864428060
        operand2 <= x"e41bdf90"; -- 3827031952
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"201c0000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fbd3b8b5"; -- 4224956597
        operand2 <= x"704bf27c"; -- 1884025468
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"50000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3b51e5ef"; -- 995223023
        operand2 <= x"e5c7cfd4"; -- 3855077332
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"5ef00000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"aa9ef683"; -- 2862544515
        operand2 <= x"6ecd742b"; -- 1858958379
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f7b41800" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9e2f8a0a"; -- 2653915658
        operand2 <= x"27cb4674"; -- 667633268
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"a0a00000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bdcfb700"; -- 3184506624
        operand2 <= x"5810dadf"; -- 1477499615
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"811933f6"; -- 2165912566
        operand2 <= x"b8ee1eaf"; -- 3102613167
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"99fb0000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0529b179"; -- 86618489
        operand2 <= x"844d37db"; -- 2219653083
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c8000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"83d942c5"; -- 2212053701
        operand2 <= x"6f10e525"; -- 1863378213
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7b2858a0" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"69d925b5"; -- 1775838645
        operand2 <= x"8ad2da70"; -- 2329074288
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"25b50000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"41f0fd1f"; -- 1106312479
        operand2 <= x"88a2350b"; -- 2292331787
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"87e8f800" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dc59cd40"; -- 3696872768
        operand2 <= x"7140493e"; -- 1900038462
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2a1d71be"; -- 706572734
        operand2 <= x"62e60ddb"; -- 1659243995
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f0000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"990a8cbc"; -- 2567605436
        operand2 <= x"7c8025e0"; -- 2088773088
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"990a8cbc" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"27a7945e"; -- 665293918
        operand2 <= x"789d6edf"; -- 2023583455
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"df7c541d"; -- 3749467165
        operand2 <= x"bc399863"; -- 3157891171
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fbe2a0e8" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"279a2984"; -- 664414596
        operand2 <= x"9228f538"; -- 2452157752
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"84000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1aab6679"; -- 447440505
        operand2 <= x"01147f2a"; -- 18120490
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ad99e400" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e3f7a57a"; -- 3824657786
        operand2 <= x"ee304c06"; -- 3996142598
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fde95e80" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c235060b"; -- 3258254859
        operand2 <= x"aff97e77"; -- 2952363639
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"05800000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f7b59017"; -- 4155871255
        operand2 <= x"84f2634e"; -- 2230477646
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6405c000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"ccb04a61"; -- 3434105441
        operand2 <= x"0b675539"; -- 191321401
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"c2000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"22524e89"; -- 575819401
        operand2 <= x"c62915bd"; -- 3324581309
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"20000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"15493ce4"; -- 357121252
        operand2 <= x"7bd10b3e"; -- 2077297470
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"153f5b6d"; -- 356473709
        operand2 <= x"5952f271"; -- 1498608241
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"b6da0000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e59615bb"; -- 3851818427
        operand2 <= x"e62e0011"; -- 3861774353
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2b760000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8563f344"; -- 2237920068
        operand2 <= x"e72d322b"; -- 3878498859
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1f9a2000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"41ee4e2b"; -- 1106136619
        operand2 <= x"2a21c544"; -- 706856260
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1ee4e2b0" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9ddad7da"; -- 2648365018
        operand2 <= x"4755da7e"; -- 1196808830
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"80000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5c1f5a28"; -- 1545558568
        operand2 <= x"38666465"; -- 946234469
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"83eb4500" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8bf9ebdf"; -- 2348411871
        operand2 <= x"9331948c"; -- 2469500044
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"9ebdf000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b125b635"; -- 2972038709
        operand2 <= x"2b414e99"; -- 725700249
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6a000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9b4c08ff"; -- 2605451519
        operand2 <= x"80d37375"; -- 2161341301
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1fe00000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c5d13947"; -- 3318823239
        operand2 <= x"6d84c403"; -- 1837417475
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"2e89ca38" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"8d39cf0f"; -- 2369376015
        operand2 <= x"ed5ba57a"; -- 3982206330
        ALUOp <= "110";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"3c000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b2278454"; -- 2988934228
        operand2 <= x"98de38f2"; -- 2564700402
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00002c89" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b2278454"; -- 2988934228
        operand2 <= x"98de38f2"; -- 2564700402
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffffec89" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"656e310c"; -- 1701720332
        operand2 <= x"b13c1618"; -- 2973505048
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000065" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"656e310c"; -- 1701720332
        operand2 <= x"b13c1618"; -- 2973505048
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000065" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a6955412"; -- 2794804242
        operand2 <= x"6c9a2dc7"; -- 1822043591
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"014d2aa8" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a6955412"; -- 2794804242
        operand2 <= x"6c9a2dc7"; -- 1822043591
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ff4d2aa8" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e429a90d"; -- 3827935501
        operand2 <= x"b8149c2f"; -- 3088358447
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0001c853" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e429a90d"; -- 3827935501
        operand2 <= x"b8149c2f"; -- 3088358447
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffffc853" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e04b812a"; -- 3763044650
        operand2 <= x"1f761506"; -- 527832326
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"03812e04" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e04b812a"; -- 3763044650
        operand2 <= x"1f761506"; -- 527832326
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ff812e04" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7edee865"; -- 2128537701
        operand2 <= x"0d8fcb47"; -- 227527495
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00fdbdd0" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7edee865"; -- 2128537701
        operand2 <= x"0d8fcb47"; -- 227527495
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00fdbdd0" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"792728f9"; -- 2032609529
        operand2 <= x"fa385126"; -- 4197994790
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"01e49ca3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"792728f9"; -- 2032609529
        operand2 <= x"fa385126"; -- 4197994790
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"01e49ca3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c1601e22"; -- 3244301858
        operand2 <= x"bda32064"; -- 3181584484
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0c1601e2" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c1601e22"; -- 3244301858
        operand2 <= x"bda32064"; -- 3181584484
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fc1601e2" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7377054b"; -- 1937179979
        operand2 <= x"a2ad9982"; -- 2729286018
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1cddc152" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7377054b"; -- 1937179979
        operand2 <= x"a2ad9982"; -- 2729286018
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1cddc152" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1267a0a9"; -- 308781225
        operand2 <= x"aba86156"; -- 2879938902
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000049" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1267a0a9"; -- 308781225
        operand2 <= x"aba86156"; -- 2879938902
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000049" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c35ffd0b"; -- 3277847819
        operand2 <= x"f3d0027c"; -- 4090495612
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000000c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c35ffd0b"; -- 3277847819
        operand2 <= x"f3d0027c"; -- 4090495612
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fffffffc" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a78bf1d0"; -- 2810966480
        operand2 <= x"11fd9161"; -- 301830497
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"53c5f8e8" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a78bf1d0"; -- 2810966480
        operand2 <= x"11fd9161"; -- 301830497
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d3c5f8e8" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7fa7f320"; -- 2141713184
        operand2 <= x"d6755b0a"; -- 3598015242
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"001fe9fc" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7fa7f320"; -- 2141713184
        operand2 <= x"d6755b0a"; -- 3598015242
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"001fe9fc" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a0f36dbb"; -- 2700307899
        operand2 <= x"5689178e"; -- 1451825038
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000283cd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"a0f36dbb"; -- 2700307899
        operand2 <= x"5689178e"; -- 1451825038
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fffe83cd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4d6bb017"; -- 1298903063
        operand2 <= x"78485260"; -- 2018005600
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4d6bb017" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4d6bb017"; -- 1298903063
        operand2 <= x"78485260"; -- 2018005600
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"4d6bb017" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"11026ea5"; -- 285372069
        operand2 <= x"da7b9252"; -- 3665531474
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000440" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"11026ea5"; -- 285372069
        operand2 <= x"da7b9252"; -- 3665531474
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000440" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"730a169f"; -- 1930040991
        operand2 <= x"a57bf93a"; -- 2776365370
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000001c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"730a169f"; -- 1930040991
        operand2 <= x"a57bf93a"; -- 2776365370
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000001c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f0c57732"; -- 4039472946
        operand2 <= x"a46ae37d"; -- 2758468477
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000007" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f0c57732"; -- 4039472946
        operand2 <= x"a46ae37d"; -- 2758468477
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffffffff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bb172756"; -- 3138856790
        operand2 <= x"45ced6fd"; -- 1171183357
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000005" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bb172756"; -- 3138856790
        operand2 <= x"45ced6fd"; -- 1171183357
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fffffffd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0c061c67"; -- 201727079
        operand2 <= x"cb1567ac"; -- 3407177644
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000c061" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0c061c67"; -- 201727079
        operand2 <= x"cb1567ac"; -- 3407177644
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000c061" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"54c758a8"; -- 1422350504
        operand2 <= x"670b48e7"; -- 1728792807
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00a98eb1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"54c758a8"; -- 1422350504
        operand2 <= x"670b48e7"; -- 1728792807
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00a98eb1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bdd1b7d8"; -- 3184637912
        operand2 <= x"f867cd8a"; -- 4167552394
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"002f746d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"bdd1b7d8"; -- 3184637912
        operand2 <= x"f867cd8a"; -- 4167552394
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffef746d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"af006d8f"; -- 2936040847
        operand2 <= x"831c9bf9"; -- 2199690233
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000057" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"af006d8f"; -- 2936040847
        operand2 <= x"831c9bf9"; -- 2199690233
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffffffd7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"eccbe6e5"; -- 3972785893
        operand2 <= x"4a22e861"; -- 1243801697
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"7665f372" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"eccbe6e5"; -- 3972785893
        operand2 <= x"4a22e861"; -- 1243801697
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f665f372" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"857d7c1a"; -- 2239593498
        operand2 <= x"aeddd388"; -- 2933773192
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00857d7c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"857d7c1a"; -- 2239593498
        operand2 <= x"aeddd388"; -- 2933773192
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ff857d7c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"acb4189b"; -- 2897483931
        operand2 <= x"53ba9301"; -- 1404736257
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"565a0c4d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"acb4189b"; -- 2897483931
        operand2 <= x"53ba9301"; -- 1404736257
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"d65a0c4d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2ec729ab"; -- 784804267
        operand2 <= x"15d2ac2a"; -- 366128170
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000bb1ca" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2ec729ab"; -- 784804267
        operand2 <= x"15d2ac2a"; -- 366128170
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000bb1ca" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"819fab35"; -- 2174724917
        operand2 <= x"8a8452a5"; -- 2323927717
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"040cfd59" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"819fab35"; -- 2174724917
        operand2 <= x"8a8452a5"; -- 2323927717
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fc0cfd59" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7a26f0e0"; -- 2049372384
        operand2 <= x"dafba573"; -- 3673924979
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000f44" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7a26f0e0"; -- 2049372384
        operand2 <= x"dafba573"; -- 3673924979
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000f44" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"19c4efb3"; -- 432336819
        operand2 <= x"4fb47ef5"; -- 1337229045
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000000ce" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"19c4efb3"; -- 432336819
        operand2 <= x"4fb47ef5"; -- 1337229045
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000000ce" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e3203449"; -- 3810538569
        operand2 <= x"b6f40274"; -- 3069444724
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000e32" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e3203449"; -- 3810538569
        operand2 <= x"b6f40274"; -- 3069444724
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fffffe32" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"da8f8579"; -- 3666838905
        operand2 <= x"eda79178"; -- 3987181944
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000000da" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"da8f8579"; -- 3666838905
        operand2 <= x"eda79178"; -- 3987181944
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffffffda" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"42f05bcf"; -- 1123048399
        operand2 <= x"5a793073"; -- 1517891699
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000085e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"42f05bcf"; -- 1123048399
        operand2 <= x"5a793073"; -- 1517891699
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000085e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0803d46f"; -- 134468719
        operand2 <= x"a5fe1f7b"; -- 2784894843
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0803d46f"; -- 134468719
        operand2 <= x"a5fe1f7b"; -- 2784894843
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1f834914"; -- 528697620
        operand2 <= x"625e2f93"; -- 1650339731
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000003f0" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1f834914"; -- 528697620
        operand2 <= x"625e2f93"; -- 1650339731
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000003f0" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d520dc15"; -- 3575700501
        operand2 <= x"f8ad1a57"; -- 4172094039
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000001aa" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d520dc15"; -- 3575700501
        operand2 <= x"f8ad1a57"; -- 4172094039
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffffffaa" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0fa71fd9"; -- 262610905
        operand2 <= x"f0b0be25"; -- 4038114853
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"007d38fe" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0fa71fd9"; -- 262610905
        operand2 <= x"f0b0be25"; -- 4038114853
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"007d38fe" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0a63920d"; -- 174297613
        operand2 <= x"7a038df9"; -- 2047053305
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000005" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0a63920d"; -- 174297613
        operand2 <= x"7a038df9"; -- 2047053305
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000005" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3210053e"; -- 839910718
        operand2 <= x"ef73202d"; -- 4017299501
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00019080" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3210053e"; -- 839910718
        operand2 <= x"ef73202d"; -- 4017299501
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00019080" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"54d38c85"; -- 1423150213
        operand2 <= x"71e74f3c"; -- 1910984508
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000005" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"54d38c85"; -- 1423150213
        operand2 <= x"71e74f3c"; -- 1910984508
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000005" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dd79b821"; -- 3715741729
        operand2 <= x"59a6e2e2"; -- 1504109282
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"375e6e08" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"dd79b821"; -- 3715741729
        operand2 <= x"59a6e2e2"; -- 1504109282
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"f75e6e08" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0c4576e8"; -- 205879016
        operand2 <= x"ea101ca9"; -- 3926924457
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000622bb" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0c4576e8"; -- 205879016
        operand2 <= x"ea101ca9"; -- 3926924457
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000622bb" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"63e4af7b"; -- 1675931515
        operand2 <= x"7780b049"; -- 2004922441
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0031f257" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"63e4af7b"; -- 1675931515
        operand2 <= x"7780b049"; -- 2004922441
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0031f257" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"61a8a9f4"; -- 1638443508
        operand2 <= x"bc6409d5"; -- 3160672725
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000030d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"61a8a9f4"; -- 1638443508
        operand2 <= x"bc6409d5"; -- 3160672725
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000030d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"841d0ecc"; -- 2216496844
        operand2 <= x"0d686918"; -- 224946456
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000084" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"841d0ecc"; -- 2216496844
        operand2 <= x"0d686918"; -- 224946456
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffffff84" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"49a11a17"; -- 1235294743
        operand2 <= x"b798615b"; -- 3080216923
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000009" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"49a11a17"; -- 1235294743
        operand2 <= x"b798615b"; -- 3080216923
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000009" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f98611a5"; -- 4186313125
        operand2 <= x"fd12f908"; -- 4245879048
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00f98611" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f98611a5"; -- 4186313125
        operand2 <= x"fd12f908"; -- 4245879048
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fff98611" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1a6dd693"; -- 443405971
        operand2 <= x"eb5556d5"; -- 3948238549
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000000d3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1a6dd693"; -- 443405971
        operand2 <= x"eb5556d5"; -- 3948238549
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000000d3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2c6afd2e"; -- 745209134
        operand2 <= x"efd38d2d"; -- 4023618861
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00016357" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2c6afd2e"; -- 745209134
        operand2 <= x"efd38d2d"; -- 4023618861
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00016357" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"26536069"; -- 642998377
        operand2 <= x"36a06239"; -- 916480569
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000013" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"26536069"; -- 642998377
        operand2 <= x"36a06239"; -- 916480569
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000013" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6524f69c"; -- 1696921244
        operand2 <= x"4746c2f3"; -- 1195819763
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000ca4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6524f69c"; -- 1696921244
        operand2 <= x"4746c2f3"; -- 1195819763
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000ca4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"18e89e96"; -- 417898134
        operand2 <= x"b9003168"; -- 3103797608
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0018e89e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"18e89e96"; -- 417898134
        operand2 <= x"b9003168"; -- 3103797608
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0018e89e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6ea6d525"; -- 1856427301
        operand2 <= x"e6a9a0b4"; -- 3869876404
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000006ea" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6ea6d525"; -- 1856427301
        operand2 <= x"e6a9a0b4"; -- 3869876404
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000006ea" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0627e208"; -- 103277064
        operand2 <= x"7ba8852d"; -- 2074641709
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000313f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0627e208"; -- 103277064
        operand2 <= x"7ba8852d"; -- 2074641709
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000313f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"effdeea0"; -- 4026396320
        operand2 <= x"52eddfae"; -- 1391321006
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0003bff7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"effdeea0"; -- 4026396320
        operand2 <= x"52eddfae"; -- 1391321006
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffffbff7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1a6b53cd"; -- 443241421
        operand2 <= x"3c717b10"; -- 1014070032
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00001a6b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1a6b53cd"; -- 443241421
        operand2 <= x"3c717b10"; -- 1014070032
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00001a6b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"28ac2c83"; -- 682372227
        operand2 <= x"e7a0bd48"; -- 3886071112
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0028ac2c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"28ac2c83"; -- 682372227
        operand2 <= x"e7a0bd48"; -- 3886071112
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0028ac2c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e5287849"; -- 3844634697
        operand2 <= x"93cb0077"; -- 2479554679
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000001ca" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e5287849"; -- 3844634697
        operand2 <= x"93cb0077"; -- 2479554679
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffffffca" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b3c16de5"; -- 3015798245
        operand2 <= x"ecd673bf"; -- 3973477311
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b3c16de5"; -- 3015798245
        operand2 <= x"ecd673bf"; -- 3973477311
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffffffff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"072d9e4f"; -- 120430159
        operand2 <= x"f273bb33"; -- 4067670835
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000000e5" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"072d9e4f"; -- 120430159
        operand2 <= x"f273bb33"; -- 4067670835
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000000e5" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e1d7f3c4"; -- 3789026244
        operand2 <= x"93c59772"; -- 2479200114
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00003875" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e1d7f3c4"; -- 3789026244
        operand2 <= x"93c59772"; -- 2479200114
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fffff875" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"30b5a59b"; -- 817210779
        operand2 <= x"7d1724e5"; -- 2098668773
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0185ad2c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"30b5a59b"; -- 817210779
        operand2 <= x"7d1724e5"; -- 2098668773
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0185ad2c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"196efc4d"; -- 426703949
        operand2 <= x"0f7de4e6"; -- 259908838
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0065bbf1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"196efc4d"; -- 426703949
        operand2 <= x"0f7de4e6"; -- 259908838
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0065bbf1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5cb6d9f7"; -- 1555487223
        operand2 <= x"52aeafcb"; -- 1387179979
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000b96db" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5cb6d9f7"; -- 1555487223
        operand2 <= x"52aeafcb"; -- 1387179979
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000b96db" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"19731df3"; -- 426974707
        operand2 <= x"f4d34250"; -- 4107485776
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00001973" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"19731df3"; -- 426974707
        operand2 <= x"f4d34250"; -- 4107485776
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00001973" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d9dda318"; -- 3655181080
        operand2 <= x"61f6b8e1"; -- 1643559137
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"6ceed18c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d9dda318"; -- 3655181080
        operand2 <= x"61f6b8e1"; -- 1643559137
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"eceed18c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b821d41c"; -- 3089224732
        operand2 <= x"7b63a768"; -- 2070128488
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00b821d4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b821d41c"; -- 3089224732
        operand2 <= x"7b63a768"; -- 2070128488
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffb821d4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7db4f3ce"; -- 2109010894
        operand2 <= x"43c5d7e3"; -- 1137039331
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0fb69e79" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7db4f3ce"; -- 2109010894
        operand2 <= x"43c5d7e3"; -- 1137039331
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0fb69e79" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"960df583"; -- 2517497219
        operand2 <= x"d913908f"; -- 3641938063
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00012c1b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"960df583"; -- 2517497219
        operand2 <= x"d913908f"; -- 3641938063
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffff2c1b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0055693f"; -- 5597503
        operand2 <= x"4bada4c6"; -- 1269671110
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000155a4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0055693f"; -- 5597503
        operand2 <= x"4bada4c6"; -- 1269671110
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000155a4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4a1c99a0"; -- 1243388320
        operand2 <= x"d4b3ec04"; -- 3568561156
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"04a1c99a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4a1c99a0"; -- 1243388320
        operand2 <= x"d4b3ec04"; -- 3568561156
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"04a1c99a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f9621693"; -- 4183955091
        operand2 <= x"92dcfa25"; -- 2463955493
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"07cb10b4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f9621693"; -- 4183955091
        operand2 <= x"92dcfa25"; -- 2463955493
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffcb10b4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"00f99a8d"; -- 16358029
        operand2 <= x"e2976736"; -- 3801573174
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000003" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"00f99a8d"; -- 16358029
        operand2 <= x"e2976736"; -- 3801573174
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000003" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"cfb7a0c4"; -- 3484917956
        operand2 <= x"7f15c8cb"; -- 2132134091
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0019f6f4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"cfb7a0c4"; -- 3484917956
        operand2 <= x"7f15c8cb"; -- 2132134091
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fff9f6f4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3b5bf67c"; -- 995882620
        operand2 <= x"7ab841fc"; -- 2058895868
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000003" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3b5bf67c"; -- 995882620
        operand2 <= x"7ab841fc"; -- 2058895868
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000003" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d0babd34"; -- 3501899060
        operand2 <= x"574747e8"; -- 1464289256
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00d0babd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d0babd34"; -- 3501899060
        operand2 <= x"574747e8"; -- 1464289256
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffd0babd" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"74c72dc5"; -- 1959210437
        operand2 <= x"048d7952"; -- 76380498
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00001d31" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"74c72dc5"; -- 1959210437
        operand2 <= x"048d7952"; -- 76380498
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00001d31" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f71a0dab"; -- 4145679787
        operand2 <= x"da2dd892"; -- 3660437650
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00003dc6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f71a0dab"; -- 4145679787
        operand2 <= x"da2dd892"; -- 3660437650
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fffffdc6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4f0e0d15"; -- 1326320917
        operand2 <= x"630486f9"; -- 1661241081
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000027" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4f0e0d15"; -- 1326320917
        operand2 <= x"630486f9"; -- 1661241081
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000027" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0a0f341d"; -- 168768541
        operand2 <= x"e4987afe"; -- 3835198206
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0a0f341d"; -- 168768541
        operand2 <= x"e4987afe"; -- 3835198206
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"eb714571"; -- 3950069105
        operand2 <= x"f00ca6c7"; -- 4027360967
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"01d6e28a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"eb714571"; -- 3950069105
        operand2 <= x"f00ca6c7"; -- 4027360967
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffd6e28a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"78e5aebe"; -- 2028318398
        operand2 <= x"641c8fcd"; -- 1679593421
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0003c72d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"78e5aebe"; -- 2028318398
        operand2 <= x"641c8fcd"; -- 1679593421
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0003c72d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"120655d7"; -- 302405079
        operand2 <= x"f09f0e5e"; -- 4036955742
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"120655d7"; -- 302405079
        operand2 <= x"f09f0e5e"; -- 4036955742
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000000" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5fde12fd"; -- 1608389373
        operand2 <= x"2209e36e"; -- 571073390
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00017f78" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5fde12fd"; -- 1608389373
        operand2 <= x"2209e36e"; -- 571073390
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00017f78" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6bdb1b93"; -- 1809521555
        operand2 <= x"da9aea35"; -- 3667585589
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000035e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6bdb1b93"; -- 1809521555
        operand2 <= x"da9aea35"; -- 3667585589
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000035e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fc31a64e"; -- 4231112270
        operand2 <= x"0872aedc"; -- 141733596
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000000f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"fc31a64e"; -- 4231112270
        operand2 <= x"0872aedc"; -- 141733596
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffffffff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b71e94d0"; -- 3072234704
        operand2 <= x"f08be826"; -- 4035700774
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"02dc7a53" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b71e94d0"; -- 3072234704
        operand2 <= x"f08be826"; -- 4035700774
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fedc7a53" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3d48c29a"; -- 1028178586
        operand2 <= x"043e4038"; -- 71188536
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000003d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3d48c29a"; -- 1028178586
        operand2 <= x"043e4038"; -- 71188536
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000003d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d9c7e253"; -- 3653755475
        operand2 <= x"db91ab79"; -- 3683756921
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000006c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d9c7e253"; -- 3653755475
        operand2 <= x"db91ab79"; -- 3683756921
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffffffec" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e3cf1286"; -- 3821998726
        operand2 <= x"d245dbc9"; -- 3527793609
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0071e789" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"e3cf1286"; -- 3821998726
        operand2 <= x"d245dbc9"; -- 3527793609
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fff1e789" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"eaaa18b1"; -- 3937015985
        operand2 <= x"89b5700b"; -- 2310369291
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"001d5543" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"eaaa18b1"; -- 3937015985
        operand2 <= x"89b5700b"; -- 2310369291
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fffd5543" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d6483feb"; -- 3595059179
        operand2 <= x"272846d9"; -- 656951001
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000006b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d6483feb"; -- 3595059179
        operand2 <= x"272846d9"; -- 656951001
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffffffeb" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1db5c0d0"; -- 498450640
        operand2 <= x"3e3af52b"; -- 1044051243
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0003b6b8" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"1db5c0d0"; -- 498450640
        operand2 <= x"3e3af52b"; -- 1044051243
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0003b6b8" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3e843304"; -- 1048851204
        operand2 <= x"9b435923"; -- 2604882211
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"07d08660" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3e843304"; -- 1048851204
        operand2 <= x"9b435923"; -- 2604882211
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"07d08660" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9bd3aaf2"; -- 2614340338
        operand2 <= x"51f3a5f0"; -- 1374922224
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00009bd3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9bd3aaf2"; -- 2614340338
        operand2 <= x"51f3a5f0"; -- 1374922224
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffff9bd3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"377665e4"; -- 930506212
        operand2 <= x"c22d894d"; -- 3257764173
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0001bbb3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"377665e4"; -- 930506212
        operand2 <= x"c22d894d"; -- 3257764173
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0001bbb3" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6e006215"; -- 1845518869
        operand2 <= x"de24fddc"; -- 3726966236
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000006" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6e006215"; -- 1845518869
        operand2 <= x"de24fddc"; -- 3726966236
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000006" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9b89d655"; -- 2609501781
        operand2 <= x"8fb849e8"; -- 2411219432
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"009b89d6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9b89d655"; -- 2609501781
        operand2 <= x"8fb849e8"; -- 2411219432
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ff9b89d6" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b440616c"; -- 3024118124
        operand2 <= x"7f355a58"; -- 2134202968
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000000b4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b440616c"; -- 3024118124
        operand2 <= x"7f355a58"; -- 2134202968
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffffffb4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9bae1293"; -- 2611876499
        operand2 <= x"7133fd4c"; -- 1899232588
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0009bae1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"9bae1293"; -- 2611876499
        operand2 <= x"7133fd4c"; -- 1899232588
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fff9bae1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"45631608"; -- 1164121608
        operand2 <= x"87973b7b"; -- 2274835323
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000008" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"45631608"; -- 1164121608
        operand2 <= x"87973b7b"; -- 2274835323
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000008" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6f64321d"; -- 1868837405
        operand2 <= x"e5ff2c1b"; -- 3858705435
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000000d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6f64321d"; -- 1868837405
        operand2 <= x"e5ff2c1b"; -- 3858705435
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000000d" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"edb279bb"; -- 3987896763
        operand2 <= x"9a3823ed"; -- 2587370477
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00076d93" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"edb279bb"; -- 3987896763
        operand2 <= x"9a3823ed"; -- 2587370477
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffff6d93" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"60fff9a1"; -- 1627388321
        operand2 <= x"e461ad23"; -- 3831606563
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0c1fff34" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"60fff9a1"; -- 1627388321
        operand2 <= x"e461ad23"; -- 3831606563
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0c1fff34" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d97477fa"; -- 3648288762
        operand2 <= x"0e2b0dd6"; -- 237702614
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000365" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"d97477fa"; -- 3648288762
        operand2 <= x"0e2b0dd6"; -- 237702614
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffffff65" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"611d50b4"; -- 1629311156
        operand2 <= x"14c4972c"; -- 348428076
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000611d5" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"611d50b4"; -- 1629311156
        operand2 <= x"14c4972c"; -- 348428076
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000611d5" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7df159dc"; -- 2112969180
        operand2 <= x"9a49337b"; -- 2588488571
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000000f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7df159dc"; -- 2112969180
        operand2 <= x"9a49337b"; -- 2588488571
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000000f" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7f0f53f1"; -- 2131710961
        operand2 <= x"a1e114a2"; -- 2715882658
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1fc3d4fc" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"7f0f53f1"; -- 2131710961
        operand2 <= x"a1e114a2"; -- 2715882658
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"1fc3d4fc" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3b50e80b"; -- 995158027
        operand2 <= x"964cd2ea"; -- 2521617130
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000ed43a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3b50e80b"; -- 995158027
        operand2 <= x"964cd2ea"; -- 2521617130
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000ed43a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5baaf8bd"; -- 1537931453
        operand2 <= x"3cced0ce"; -- 1020186830
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00016eab" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"5baaf8bd"; -- 1537931453
        operand2 <= x"3cced0ce"; -- 1020186830
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00016eab" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3be68ce8"; -- 1004965096
        operand2 <= x"f78fe9bc"; -- 4153403836
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000003" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3be68ce8"; -- 1004965096
        operand2 <= x"f78fe9bc"; -- 4153403836
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000003" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"570bbe24"; -- 1460387364
        operand2 <= x"6f9ca4ce"; -- 1872536782
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00015c2e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"570bbe24"; -- 1460387364
        operand2 <= x"6f9ca4ce"; -- 1872536782
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00015c2e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6b52758f"; -- 1800566159
        operand2 <= x"b22f03a3"; -- 2989425571
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0d6a4eb1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"6b52758f"; -- 1800566159
        operand2 <= x"b22f03a3"; -- 2989425571
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0d6a4eb1" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"42000380"; -- 1107297152
        operand2 <= x"d9a98c75"; -- 3651767413
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000210" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"42000380"; -- 1107297152
        operand2 <= x"d9a98c75"; -- 3651767413
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000210" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4494374f"; -- 1150564175
        operand2 <= x"31f13823"; -- 837892131
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"089286e9" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"4494374f"; -- 1150564175
        operand2 <= x"31f13823"; -- 837892131
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"089286e9" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f961ad0a"; -- 4183928074
        operand2 <= x"82259606"; -- 2183501318
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"03e586b4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"f961ad0a"; -- 4183928074
        operand2 <= x"82259606"; -- 2183501318
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffe586b4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"614f5722"; -- 1632589602
        operand2 <= x"4799330d"; -- 1201222413
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00030a7a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"614f5722"; -- 1632589602
        operand2 <= x"4799330d"; -- 1201222413
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00030a7a" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b941be17"; -- 3108093463
        operand2 <= x"99f16029"; -- 2582732841
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"005ca0df" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b941be17"; -- 3108093463
        operand2 <= x"99f16029"; -- 2582732841
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffdca0df" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c5df8dad"; -- 3319762349
        operand2 <= x"e737a635"; -- 3879183925
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000062e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"c5df8dad"; -- 3319762349
        operand2 <= x"e737a635"; -- 3879183925
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"fffffe2e" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"18d8bbef"; -- 416857071
        operand2 <= x"2d6da28c"; -- 762159756
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00018d8b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"18d8bbef"; -- 416857071
        operand2 <= x"2d6da28c"; -- 762159756
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00018d8b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3b53d175"; -- 995348853
        operand2 <= x"5959040a"; -- 1499005962
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000ed4f4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"3b53d175"; -- 995348853
        operand2 <= x"5959040a"; -- 1499005962
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000ed4f4" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2d89ef95"; -- 764014485
        operand2 <= x"3f52354a"; -- 1062352202
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000b627b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"2d89ef95"; -- 764014485
        operand2 <= x"3f52354a"; -- 1062352202
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"000b627b" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b9ce97b4"; -- 3117324212
        operand2 <= x"982e261f"; -- 2553161247
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00000001" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"b9ce97b4"; -- 3117324212
        operand2 <= x"982e261f"; -- 2553161247
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"ffffffff" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"47fafe5b"; -- 1207631451
        operand2 <= x"49ed31cd"; -- 1240281549
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00023fd7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"47fafe5b"; -- 1207631451
        operand2 <= x"49ed31cd"; -- 1240281549
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"00023fd7" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0c572d28"; -- 207039784
        operand2 <= x"6f2f84f8"; -- 1865385208
        ALUOp <= "111";
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000000c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        -- apply stimuli
        operand1 <= x"0c572d28"; -- 207039784
        operand2 <= x"6f2f84f8"; -- 1865385208
        ALUOp <= "111";
        arith_logic_b <= '1';
        signed_unsigned_b <= '0';
        wait for 2 ns;
        -- check outputs
        if result /= x"0000000c" then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if equal /= '0' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_u /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        if x_lt_y_s /= '1' then
            bad_checks := bad_checks + 1;
        else
            good_checks := good_checks + 1;
        end if;
        wait for 2 ns;

        operand1 <= (others => '0');
        operand2 <= (others => '0');
        ALUOp <= (others => '0');
        arith_logic_b <= '0';
        signed_unsigned_b <= '0';
        report "DISCH_GRADING (good, bad, total): " & integer'image(good_checks) & " " & integer'image(bad_checks) & " " & integer'image(good_checks + bad_checks) & "" severity note;

        wait;
    end process;

    DUT: component alu port map(
        operand1 => operand1,
        operand2 => operand2,
        ALUOp => ALUOp,
        arith_logic_b => arith_logic_b,
        signed_unsigned_b => signed_unsigned_b,
        result => result,
        equal => equal,
        x_lt_y_u => x_lt_y_u,
        x_lt_y_s => x_lt_y_s
    );

end Behavioural;
